magic
tech sky130A
magscale 1 2
timestamp 1741017040
<< viali >>
rect 43361 101609 43395 101643
rect 45293 101609 45327 101643
rect 47961 101609 47995 101643
rect 49893 101609 49927 101643
rect 51089 101609 51123 101643
rect 53021 101609 53055 101643
rect 55689 101609 55723 101643
rect 57621 101609 57655 101643
rect 58817 101609 58851 101643
rect 43545 101405 43579 101439
rect 45477 101405 45511 101439
rect 47777 101405 47811 101439
rect 49709 101405 49743 101439
rect 51273 101405 51307 101439
rect 53205 101405 53239 101439
rect 55505 101405 55539 101439
rect 57437 101405 57471 101439
rect 59001 101405 59035 101439
rect 43545 77673 43579 77707
rect 47501 77673 47535 77707
rect 49709 77673 49743 77707
rect 53113 77673 53147 77707
rect 55137 77673 55171 77707
rect 57345 77673 57379 77707
rect 59185 77673 59219 77707
rect 41797 77537 41831 77571
rect 45753 77537 45787 77571
rect 47961 77537 47995 77571
rect 51365 77537 51399 77571
rect 53389 77537 53423 77571
rect 55597 77537 55631 77571
rect 57437 77537 57471 77571
rect 42073 77401 42107 77435
rect 46029 77401 46063 77435
rect 48237 77401 48271 77435
rect 51641 77401 51675 77435
rect 53665 77401 53699 77435
rect 55873 77401 55907 77435
rect 57713 77401 57747 77435
rect 41705 77333 41739 77367
rect 45385 77129 45419 77163
rect 51181 77129 51215 77163
rect 49709 77061 49743 77095
rect 43637 76993 43671 77027
rect 49433 76993 49467 77027
rect 43913 76925 43947 76959
rect 41797 76789 41831 76823
rect 45753 76789 45787 76823
rect 47961 76789 47995 76823
rect 51365 76789 51399 76823
rect 53389 76789 53423 76823
rect 55597 76789 55631 76823
rect 57529 76789 57563 76823
rect 49525 76585 49559 76619
rect 43637 76245 43671 76279
rect 46581 74953 46615 74987
rect 48237 74953 48271 74987
rect 49985 74953 50019 74987
rect 51917 74953 51951 74987
rect 53205 74953 53239 74987
rect 54861 74953 54895 74987
rect 56885 74953 56919 74987
rect 58357 74953 58391 74987
rect 60657 74953 60691 74987
rect 46673 74817 46707 74851
rect 48329 74817 48363 74851
rect 50077 74817 50111 74851
rect 52009 74817 52043 74851
rect 53297 74817 53331 74851
rect 54953 74817 54987 74851
rect 56977 74817 57011 74851
rect 58449 74817 58483 74851
rect 60197 74817 60231 74851
rect 60473 74817 60507 74851
rect 60565 74817 60599 74851
rect 100217 62849 100251 62883
rect 100401 62645 100435 62679
rect 1685 62237 1719 62271
rect 100217 62237 100251 62271
rect 1501 62101 1535 62135
rect 1869 62101 1903 62135
rect 100401 62101 100435 62135
rect 1685 61761 1719 61795
rect 100217 61761 100251 61795
rect 1501 61557 1535 61591
rect 100401 61557 100435 61591
rect 21097 61353 21131 61387
rect 81909 61353 81943 61387
rect 82350 61353 82384 61387
rect 22569 61217 22603 61251
rect 78873 61217 78907 61251
rect 80621 61217 80655 61251
rect 22845 61149 22879 61183
rect 77033 61149 77067 61183
rect 80713 61149 80747 61183
rect 82093 61149 82127 61183
rect 83933 61149 83967 61183
rect 77309 61081 77343 61115
rect 79149 61081 79183 61115
rect 76849 61013 76883 61047
rect 78781 61013 78815 61047
rect 83841 61013 83875 61047
rect 84025 61013 84059 61047
rect 30389 60809 30423 60843
rect 48145 60741 48179 60775
rect 29193 60673 29227 60707
rect 29285 60673 29319 60707
rect 30481 60673 30515 60707
rect 77217 60673 77251 60707
rect 78505 60673 78539 60707
rect 79241 60673 79275 60707
rect 79333 60673 79367 60707
rect 79701 60673 79735 60707
rect 100217 60673 100251 60707
rect 24041 60605 24075 60639
rect 24317 60605 24351 60639
rect 77125 60605 77159 60639
rect 78597 60605 78631 60639
rect 79977 60605 80011 60639
rect 81541 60605 81575 60639
rect 81817 60605 81851 60639
rect 83381 60605 83415 60639
rect 83933 60605 83967 60639
rect 85681 60605 85715 60639
rect 85957 60605 85991 60639
rect 87613 60605 87647 60639
rect 87889 60605 87923 60639
rect 22569 60537 22603 60571
rect 100401 60537 100435 60571
rect 22385 60469 22419 60503
rect 79517 60469 79551 60503
rect 81449 60469 81483 60503
rect 83289 60469 83323 60503
rect 86141 60469 86175 60503
rect 48421 60265 48455 60299
rect 80253 60265 80287 60299
rect 81817 60265 81851 60299
rect 84485 60265 84519 60299
rect 85957 60265 85991 60299
rect 87705 60265 87739 60299
rect 75469 60129 75503 60163
rect 85129 60129 85163 60163
rect 87613 60129 87647 60163
rect 87981 60129 88015 60163
rect 80161 60061 80195 60095
rect 81725 60061 81759 60095
rect 84393 60061 84427 60095
rect 85773 60061 85807 60095
rect 85865 60061 85899 60095
rect 86969 60061 87003 60095
rect 88073 60061 88107 60095
rect 100217 60061 100251 60095
rect 49893 59993 49927 60027
rect 57069 59993 57103 60027
rect 73721 59993 73755 60027
rect 55781 59925 55815 59959
rect 100401 59925 100435 59959
rect 98285 53941 98319 53975
rect 98561 46053 98595 46087
rect 98285 45917 98319 45951
rect 98377 45917 98411 45951
rect 98561 45849 98595 45883
rect 98469 45033 98503 45067
rect 98285 44761 98319 44795
rect 98469 44693 98503 44727
rect 98653 44693 98687 44727
rect 98285 43265 98319 43299
rect 98377 43061 98411 43095
rect 99849 41021 99883 41055
rect 100125 41021 100159 41055
rect 98377 40885 98411 40919
rect 98469 40681 98503 40715
rect 98285 40477 98319 40511
rect 98469 40477 98503 40511
rect 98285 35649 98319 35683
rect 98377 35445 98411 35479
rect 98285 34561 98319 34595
rect 98377 34493 98411 34527
rect 98377 31841 98411 31875
rect 99849 31841 99883 31875
rect 100125 31773 100159 31807
rect 100033 30685 100067 30719
rect 99757 30617 99791 30651
rect 98285 30549 98319 30583
rect 98837 30209 98871 30243
rect 99389 30005 99423 30039
rect 98285 29597 98319 29631
rect 98377 29461 98411 29495
rect 98377 29121 98411 29155
rect 99941 29121 99975 29155
rect 98929 29053 98963 29087
rect 99849 29053 99883 29087
rect 98469 28985 98503 29019
rect 99481 28985 99515 29019
rect 99573 28985 99607 29019
rect 99665 27557 99699 27591
rect 99389 27489 99423 27523
rect 99849 27489 99883 27523
rect 99297 27421 99331 27455
rect 99757 27421 99791 27455
rect 99941 27421 99975 27455
rect 100309 26469 100343 26503
rect 98653 26401 98687 26435
rect 98929 26333 98963 26367
rect 100493 26333 100527 26367
rect 99552 25993 99586 26027
rect 98377 25925 98411 25959
rect 99757 25925 99791 25959
rect 99113 25789 99147 25823
rect 99389 25653 99423 25687
rect 99573 25653 99607 25687
rect 99849 25313 99883 25347
rect 100125 25245 100159 25279
rect 98377 25109 98411 25143
rect 99941 24701 99975 24735
rect 100217 24701 100251 24735
rect 98469 24565 98503 24599
rect 98377 24157 98411 24191
rect 98469 24021 98503 24055
rect 98745 23817 98779 23851
rect 98929 23817 98963 23851
rect 98285 23681 98319 23715
rect 98804 23681 98838 23715
rect 98377 23477 98411 23511
rect 98485 22729 98519 22763
rect 98653 22729 98687 22763
rect 99389 22729 99423 22763
rect 98285 22661 98319 22695
rect 98837 22661 98871 22695
rect 98745 22593 98779 22627
rect 99021 22593 99055 22627
rect 99297 22593 99331 22627
rect 99481 22593 99515 22627
rect 99021 22457 99055 22491
rect 98469 22389 98503 22423
rect 98469 22185 98503 22219
rect 98285 21913 98319 21947
rect 98501 21913 98535 21947
rect 98653 21845 98687 21879
rect 99849 19873 99883 19907
rect 100125 19873 100159 19907
rect 98377 19669 98411 19703
rect 99021 19261 99055 19295
rect 98469 19125 98503 19159
rect 98469 18241 98503 18275
rect 98561 18173 98595 18207
rect 98837 18173 98871 18207
<< metal1 >>
rect 1104 101754 100832 101776
rect 1104 101702 4214 101754
rect 4266 101702 4278 101754
rect 4330 101702 4342 101754
rect 4394 101702 4406 101754
rect 4458 101702 4470 101754
rect 4522 101702 34934 101754
rect 34986 101702 34998 101754
rect 35050 101702 35062 101754
rect 35114 101702 35126 101754
rect 35178 101702 35190 101754
rect 35242 101702 65654 101754
rect 65706 101702 65718 101754
rect 65770 101702 65782 101754
rect 65834 101702 65846 101754
rect 65898 101702 65910 101754
rect 65962 101702 96374 101754
rect 96426 101702 96438 101754
rect 96490 101702 96502 101754
rect 96554 101702 96566 101754
rect 96618 101702 96630 101754
rect 96682 101702 100832 101754
rect 1104 101680 100832 101702
rect 43346 101600 43352 101652
rect 43404 101600 43410 101652
rect 45278 101600 45284 101652
rect 45336 101600 45342 101652
rect 47946 101600 47952 101652
rect 48004 101600 48010 101652
rect 49510 101600 49516 101652
rect 49568 101640 49574 101652
rect 49881 101643 49939 101649
rect 49881 101640 49893 101643
rect 49568 101612 49893 101640
rect 49568 101600 49574 101612
rect 49881 101609 49893 101612
rect 49927 101609 49939 101643
rect 49881 101603 49939 101609
rect 50982 101600 50988 101652
rect 51040 101640 51046 101652
rect 51077 101643 51135 101649
rect 51077 101640 51089 101643
rect 51040 101612 51089 101640
rect 51040 101600 51046 101612
rect 51077 101609 51089 101612
rect 51123 101609 51135 101643
rect 51077 101603 51135 101609
rect 53006 101600 53012 101652
rect 53064 101600 53070 101652
rect 55674 101600 55680 101652
rect 55732 101600 55738 101652
rect 57606 101600 57612 101652
rect 57664 101600 57670 101652
rect 58802 101600 58808 101652
rect 58860 101600 58866 101652
rect 43530 101396 43536 101448
rect 43588 101396 43594 101448
rect 45370 101396 45376 101448
rect 45428 101436 45434 101448
rect 45465 101439 45523 101445
rect 45465 101436 45477 101439
rect 45428 101408 45477 101436
rect 45428 101396 45434 101408
rect 45465 101405 45477 101408
rect 45511 101405 45523 101439
rect 45465 101399 45523 101405
rect 47486 101396 47492 101448
rect 47544 101436 47550 101448
rect 47765 101439 47823 101445
rect 47765 101436 47777 101439
rect 47544 101408 47777 101436
rect 47544 101396 47550 101408
rect 47765 101405 47777 101408
rect 47811 101405 47823 101439
rect 47765 101399 47823 101405
rect 49694 101396 49700 101448
rect 49752 101396 49758 101448
rect 51166 101396 51172 101448
rect 51224 101436 51230 101448
rect 51261 101439 51319 101445
rect 51261 101436 51273 101439
rect 51224 101408 51273 101436
rect 51224 101396 51230 101408
rect 51261 101405 51273 101408
rect 51307 101405 51319 101439
rect 51261 101399 51319 101405
rect 53098 101396 53104 101448
rect 53156 101436 53162 101448
rect 53193 101439 53251 101445
rect 53193 101436 53205 101439
rect 53156 101408 53205 101436
rect 53156 101396 53162 101408
rect 53193 101405 53205 101408
rect 53239 101405 53251 101439
rect 53193 101399 53251 101405
rect 55122 101396 55128 101448
rect 55180 101436 55186 101448
rect 55493 101439 55551 101445
rect 55493 101436 55505 101439
rect 55180 101408 55505 101436
rect 55180 101396 55186 101408
rect 55493 101405 55505 101408
rect 55539 101405 55551 101439
rect 55493 101399 55551 101405
rect 57330 101396 57336 101448
rect 57388 101436 57394 101448
rect 57425 101439 57483 101445
rect 57425 101436 57437 101439
rect 57388 101408 57437 101436
rect 57388 101396 57394 101408
rect 57425 101405 57437 101408
rect 57471 101405 57483 101439
rect 57425 101399 57483 101405
rect 58989 101439 59047 101445
rect 58989 101405 59001 101439
rect 59035 101436 59047 101439
rect 59170 101436 59176 101448
rect 59035 101408 59176 101436
rect 59035 101405 59047 101408
rect 58989 101399 59047 101405
rect 59170 101396 59176 101408
rect 59228 101396 59234 101448
rect 1104 101210 100832 101232
rect 1104 101158 4874 101210
rect 4926 101158 4938 101210
rect 4990 101158 5002 101210
rect 5054 101158 5066 101210
rect 5118 101158 5130 101210
rect 5182 101158 35594 101210
rect 35646 101158 35658 101210
rect 35710 101158 35722 101210
rect 35774 101158 35786 101210
rect 35838 101158 35850 101210
rect 35902 101158 66314 101210
rect 66366 101158 66378 101210
rect 66430 101158 66442 101210
rect 66494 101158 66506 101210
rect 66558 101158 66570 101210
rect 66622 101158 97034 101210
rect 97086 101158 97098 101210
rect 97150 101158 97162 101210
rect 97214 101158 97226 101210
rect 97278 101158 97290 101210
rect 97342 101158 100832 101210
rect 1104 101136 100832 101158
rect 1104 100666 100832 100688
rect 1104 100614 4214 100666
rect 4266 100614 4278 100666
rect 4330 100614 4342 100666
rect 4394 100614 4406 100666
rect 4458 100614 4470 100666
rect 4522 100614 34934 100666
rect 34986 100614 34998 100666
rect 35050 100614 35062 100666
rect 35114 100614 35126 100666
rect 35178 100614 35190 100666
rect 35242 100614 65654 100666
rect 65706 100614 65718 100666
rect 65770 100614 65782 100666
rect 65834 100614 65846 100666
rect 65898 100614 65910 100666
rect 65962 100614 96374 100666
rect 96426 100614 96438 100666
rect 96490 100614 96502 100666
rect 96554 100614 96566 100666
rect 96618 100614 96630 100666
rect 96682 100614 100832 100666
rect 1104 100592 100832 100614
rect 1104 100122 100832 100144
rect 1104 100070 4874 100122
rect 4926 100070 4938 100122
rect 4990 100070 5002 100122
rect 5054 100070 5066 100122
rect 5118 100070 5130 100122
rect 5182 100070 35594 100122
rect 35646 100070 35658 100122
rect 35710 100070 35722 100122
rect 35774 100070 35786 100122
rect 35838 100070 35850 100122
rect 35902 100070 66314 100122
rect 66366 100070 66378 100122
rect 66430 100070 66442 100122
rect 66494 100070 66506 100122
rect 66558 100070 66570 100122
rect 66622 100070 97034 100122
rect 97086 100070 97098 100122
rect 97150 100070 97162 100122
rect 97214 100070 97226 100122
rect 97278 100070 97290 100122
rect 97342 100070 100832 100122
rect 1104 100048 100832 100070
rect 1104 99578 100832 99600
rect 1104 99526 4214 99578
rect 4266 99526 4278 99578
rect 4330 99526 4342 99578
rect 4394 99526 4406 99578
rect 4458 99526 4470 99578
rect 4522 99526 34934 99578
rect 34986 99526 34998 99578
rect 35050 99526 35062 99578
rect 35114 99526 35126 99578
rect 35178 99526 35190 99578
rect 35242 99526 65654 99578
rect 65706 99526 65718 99578
rect 65770 99526 65782 99578
rect 65834 99526 65846 99578
rect 65898 99526 65910 99578
rect 65962 99526 96374 99578
rect 96426 99526 96438 99578
rect 96490 99526 96502 99578
rect 96554 99526 96566 99578
rect 96618 99526 96630 99578
rect 96682 99526 100832 99578
rect 1104 99504 100832 99526
rect 1104 99034 100832 99056
rect 1104 98982 4874 99034
rect 4926 98982 4938 99034
rect 4990 98982 5002 99034
rect 5054 98982 5066 99034
rect 5118 98982 5130 99034
rect 5182 98982 35594 99034
rect 35646 98982 35658 99034
rect 35710 98982 35722 99034
rect 35774 98982 35786 99034
rect 35838 98982 35850 99034
rect 35902 98982 66314 99034
rect 66366 98982 66378 99034
rect 66430 98982 66442 99034
rect 66494 98982 66506 99034
rect 66558 98982 66570 99034
rect 66622 98982 97034 99034
rect 97086 98982 97098 99034
rect 97150 98982 97162 99034
rect 97214 98982 97226 99034
rect 97278 98982 97290 99034
rect 97342 98982 100832 99034
rect 1104 98960 100832 98982
rect 1104 98490 100832 98512
rect 1104 98438 4214 98490
rect 4266 98438 4278 98490
rect 4330 98438 4342 98490
rect 4394 98438 4406 98490
rect 4458 98438 4470 98490
rect 4522 98438 34934 98490
rect 34986 98438 34998 98490
rect 35050 98438 35062 98490
rect 35114 98438 35126 98490
rect 35178 98438 35190 98490
rect 35242 98438 65654 98490
rect 65706 98438 65718 98490
rect 65770 98438 65782 98490
rect 65834 98438 65846 98490
rect 65898 98438 65910 98490
rect 65962 98438 96374 98490
rect 96426 98438 96438 98490
rect 96490 98438 96502 98490
rect 96554 98438 96566 98490
rect 96618 98438 96630 98490
rect 96682 98438 100832 98490
rect 1104 98416 100832 98438
rect 1104 97946 100832 97968
rect 1104 97894 4874 97946
rect 4926 97894 4938 97946
rect 4990 97894 5002 97946
rect 5054 97894 5066 97946
rect 5118 97894 5130 97946
rect 5182 97894 35594 97946
rect 35646 97894 35658 97946
rect 35710 97894 35722 97946
rect 35774 97894 35786 97946
rect 35838 97894 35850 97946
rect 35902 97894 66314 97946
rect 66366 97894 66378 97946
rect 66430 97894 66442 97946
rect 66494 97894 66506 97946
rect 66558 97894 66570 97946
rect 66622 97894 97034 97946
rect 97086 97894 97098 97946
rect 97150 97894 97162 97946
rect 97214 97894 97226 97946
rect 97278 97894 97290 97946
rect 97342 97894 100832 97946
rect 1104 97872 100832 97894
rect 1104 97402 100832 97424
rect 1104 97350 4214 97402
rect 4266 97350 4278 97402
rect 4330 97350 4342 97402
rect 4394 97350 4406 97402
rect 4458 97350 4470 97402
rect 4522 97350 34934 97402
rect 34986 97350 34998 97402
rect 35050 97350 35062 97402
rect 35114 97350 35126 97402
rect 35178 97350 35190 97402
rect 35242 97350 65654 97402
rect 65706 97350 65718 97402
rect 65770 97350 65782 97402
rect 65834 97350 65846 97402
rect 65898 97350 65910 97402
rect 65962 97350 96374 97402
rect 96426 97350 96438 97402
rect 96490 97350 96502 97402
rect 96554 97350 96566 97402
rect 96618 97350 96630 97402
rect 96682 97350 100832 97402
rect 1104 97328 100832 97350
rect 1104 96858 100832 96880
rect 1104 96806 4874 96858
rect 4926 96806 4938 96858
rect 4990 96806 5002 96858
rect 5054 96806 5066 96858
rect 5118 96806 5130 96858
rect 5182 96806 35594 96858
rect 35646 96806 35658 96858
rect 35710 96806 35722 96858
rect 35774 96806 35786 96858
rect 35838 96806 35850 96858
rect 35902 96806 66314 96858
rect 66366 96806 66378 96858
rect 66430 96806 66442 96858
rect 66494 96806 66506 96858
rect 66558 96806 66570 96858
rect 66622 96806 97034 96858
rect 97086 96806 97098 96858
rect 97150 96806 97162 96858
rect 97214 96806 97226 96858
rect 97278 96806 97290 96858
rect 97342 96806 100832 96858
rect 1104 96784 100832 96806
rect 1104 96314 100832 96336
rect 1104 96262 4214 96314
rect 4266 96262 4278 96314
rect 4330 96262 4342 96314
rect 4394 96262 4406 96314
rect 4458 96262 4470 96314
rect 4522 96262 34934 96314
rect 34986 96262 34998 96314
rect 35050 96262 35062 96314
rect 35114 96262 35126 96314
rect 35178 96262 35190 96314
rect 35242 96262 65654 96314
rect 65706 96262 65718 96314
rect 65770 96262 65782 96314
rect 65834 96262 65846 96314
rect 65898 96262 65910 96314
rect 65962 96262 96374 96314
rect 96426 96262 96438 96314
rect 96490 96262 96502 96314
rect 96554 96262 96566 96314
rect 96618 96262 96630 96314
rect 96682 96262 100832 96314
rect 1104 96240 100832 96262
rect 1104 95770 100832 95792
rect 1104 95718 4874 95770
rect 4926 95718 4938 95770
rect 4990 95718 5002 95770
rect 5054 95718 5066 95770
rect 5118 95718 5130 95770
rect 5182 95718 35594 95770
rect 35646 95718 35658 95770
rect 35710 95718 35722 95770
rect 35774 95718 35786 95770
rect 35838 95718 35850 95770
rect 35902 95718 66314 95770
rect 66366 95718 66378 95770
rect 66430 95718 66442 95770
rect 66494 95718 66506 95770
rect 66558 95718 66570 95770
rect 66622 95718 97034 95770
rect 97086 95718 97098 95770
rect 97150 95718 97162 95770
rect 97214 95718 97226 95770
rect 97278 95718 97290 95770
rect 97342 95718 100832 95770
rect 1104 95696 100832 95718
rect 1104 95226 100832 95248
rect 1104 95174 4214 95226
rect 4266 95174 4278 95226
rect 4330 95174 4342 95226
rect 4394 95174 4406 95226
rect 4458 95174 4470 95226
rect 4522 95174 34934 95226
rect 34986 95174 34998 95226
rect 35050 95174 35062 95226
rect 35114 95174 35126 95226
rect 35178 95174 35190 95226
rect 35242 95174 65654 95226
rect 65706 95174 65718 95226
rect 65770 95174 65782 95226
rect 65834 95174 65846 95226
rect 65898 95174 65910 95226
rect 65962 95174 96374 95226
rect 96426 95174 96438 95226
rect 96490 95174 96502 95226
rect 96554 95174 96566 95226
rect 96618 95174 96630 95226
rect 96682 95174 100832 95226
rect 1104 95152 100832 95174
rect 1104 94682 100832 94704
rect 1104 94630 4874 94682
rect 4926 94630 4938 94682
rect 4990 94630 5002 94682
rect 5054 94630 5066 94682
rect 5118 94630 5130 94682
rect 5182 94630 35594 94682
rect 35646 94630 35658 94682
rect 35710 94630 35722 94682
rect 35774 94630 35786 94682
rect 35838 94630 35850 94682
rect 35902 94630 66314 94682
rect 66366 94630 66378 94682
rect 66430 94630 66442 94682
rect 66494 94630 66506 94682
rect 66558 94630 66570 94682
rect 66622 94630 97034 94682
rect 97086 94630 97098 94682
rect 97150 94630 97162 94682
rect 97214 94630 97226 94682
rect 97278 94630 97290 94682
rect 97342 94630 100832 94682
rect 1104 94608 100832 94630
rect 1104 94138 100832 94160
rect 1104 94086 4214 94138
rect 4266 94086 4278 94138
rect 4330 94086 4342 94138
rect 4394 94086 4406 94138
rect 4458 94086 4470 94138
rect 4522 94086 34934 94138
rect 34986 94086 34998 94138
rect 35050 94086 35062 94138
rect 35114 94086 35126 94138
rect 35178 94086 35190 94138
rect 35242 94086 65654 94138
rect 65706 94086 65718 94138
rect 65770 94086 65782 94138
rect 65834 94086 65846 94138
rect 65898 94086 65910 94138
rect 65962 94086 96374 94138
rect 96426 94086 96438 94138
rect 96490 94086 96502 94138
rect 96554 94086 96566 94138
rect 96618 94086 96630 94138
rect 96682 94086 100832 94138
rect 1104 94064 100832 94086
rect 1104 93594 100832 93616
rect 1104 93542 4874 93594
rect 4926 93542 4938 93594
rect 4990 93542 5002 93594
rect 5054 93542 5066 93594
rect 5118 93542 5130 93594
rect 5182 93542 35594 93594
rect 35646 93542 35658 93594
rect 35710 93542 35722 93594
rect 35774 93542 35786 93594
rect 35838 93542 35850 93594
rect 35902 93542 66314 93594
rect 66366 93542 66378 93594
rect 66430 93542 66442 93594
rect 66494 93542 66506 93594
rect 66558 93542 66570 93594
rect 66622 93542 97034 93594
rect 97086 93542 97098 93594
rect 97150 93542 97162 93594
rect 97214 93542 97226 93594
rect 97278 93542 97290 93594
rect 97342 93542 100832 93594
rect 1104 93520 100832 93542
rect 1104 93050 100832 93072
rect 1104 92998 4214 93050
rect 4266 92998 4278 93050
rect 4330 92998 4342 93050
rect 4394 92998 4406 93050
rect 4458 92998 4470 93050
rect 4522 92998 34934 93050
rect 34986 92998 34998 93050
rect 35050 92998 35062 93050
rect 35114 92998 35126 93050
rect 35178 92998 35190 93050
rect 35242 92998 65654 93050
rect 65706 92998 65718 93050
rect 65770 92998 65782 93050
rect 65834 92998 65846 93050
rect 65898 92998 65910 93050
rect 65962 92998 96374 93050
rect 96426 92998 96438 93050
rect 96490 92998 96502 93050
rect 96554 92998 96566 93050
rect 96618 92998 96630 93050
rect 96682 92998 100832 93050
rect 1104 92976 100832 92998
rect 1104 92506 100832 92528
rect 1104 92454 4874 92506
rect 4926 92454 4938 92506
rect 4990 92454 5002 92506
rect 5054 92454 5066 92506
rect 5118 92454 5130 92506
rect 5182 92454 35594 92506
rect 35646 92454 35658 92506
rect 35710 92454 35722 92506
rect 35774 92454 35786 92506
rect 35838 92454 35850 92506
rect 35902 92454 66314 92506
rect 66366 92454 66378 92506
rect 66430 92454 66442 92506
rect 66494 92454 66506 92506
rect 66558 92454 66570 92506
rect 66622 92454 97034 92506
rect 97086 92454 97098 92506
rect 97150 92454 97162 92506
rect 97214 92454 97226 92506
rect 97278 92454 97290 92506
rect 97342 92454 100832 92506
rect 1104 92432 100832 92454
rect 1104 91962 100832 91984
rect 1104 91910 4214 91962
rect 4266 91910 4278 91962
rect 4330 91910 4342 91962
rect 4394 91910 4406 91962
rect 4458 91910 4470 91962
rect 4522 91910 34934 91962
rect 34986 91910 34998 91962
rect 35050 91910 35062 91962
rect 35114 91910 35126 91962
rect 35178 91910 35190 91962
rect 35242 91910 65654 91962
rect 65706 91910 65718 91962
rect 65770 91910 65782 91962
rect 65834 91910 65846 91962
rect 65898 91910 65910 91962
rect 65962 91910 96374 91962
rect 96426 91910 96438 91962
rect 96490 91910 96502 91962
rect 96554 91910 96566 91962
rect 96618 91910 96630 91962
rect 96682 91910 100832 91962
rect 1104 91888 100832 91910
rect 1104 91418 100832 91440
rect 1104 91366 4874 91418
rect 4926 91366 4938 91418
rect 4990 91366 5002 91418
rect 5054 91366 5066 91418
rect 5118 91366 5130 91418
rect 5182 91366 35594 91418
rect 35646 91366 35658 91418
rect 35710 91366 35722 91418
rect 35774 91366 35786 91418
rect 35838 91366 35850 91418
rect 35902 91366 66314 91418
rect 66366 91366 66378 91418
rect 66430 91366 66442 91418
rect 66494 91366 66506 91418
rect 66558 91366 66570 91418
rect 66622 91366 97034 91418
rect 97086 91366 97098 91418
rect 97150 91366 97162 91418
rect 97214 91366 97226 91418
rect 97278 91366 97290 91418
rect 97342 91366 100832 91418
rect 1104 91344 100832 91366
rect 1104 90874 100832 90896
rect 1104 90822 4214 90874
rect 4266 90822 4278 90874
rect 4330 90822 4342 90874
rect 4394 90822 4406 90874
rect 4458 90822 4470 90874
rect 4522 90822 34934 90874
rect 34986 90822 34998 90874
rect 35050 90822 35062 90874
rect 35114 90822 35126 90874
rect 35178 90822 35190 90874
rect 35242 90822 65654 90874
rect 65706 90822 65718 90874
rect 65770 90822 65782 90874
rect 65834 90822 65846 90874
rect 65898 90822 65910 90874
rect 65962 90822 96374 90874
rect 96426 90822 96438 90874
rect 96490 90822 96502 90874
rect 96554 90822 96566 90874
rect 96618 90822 96630 90874
rect 96682 90822 100832 90874
rect 1104 90800 100832 90822
rect 1104 90330 100832 90352
rect 1104 90278 4874 90330
rect 4926 90278 4938 90330
rect 4990 90278 5002 90330
rect 5054 90278 5066 90330
rect 5118 90278 5130 90330
rect 5182 90278 35594 90330
rect 35646 90278 35658 90330
rect 35710 90278 35722 90330
rect 35774 90278 35786 90330
rect 35838 90278 35850 90330
rect 35902 90278 66314 90330
rect 66366 90278 66378 90330
rect 66430 90278 66442 90330
rect 66494 90278 66506 90330
rect 66558 90278 66570 90330
rect 66622 90278 97034 90330
rect 97086 90278 97098 90330
rect 97150 90278 97162 90330
rect 97214 90278 97226 90330
rect 97278 90278 97290 90330
rect 97342 90278 100832 90330
rect 1104 90256 100832 90278
rect 1104 89786 100832 89808
rect 1104 89734 4214 89786
rect 4266 89734 4278 89786
rect 4330 89734 4342 89786
rect 4394 89734 4406 89786
rect 4458 89734 4470 89786
rect 4522 89734 34934 89786
rect 34986 89734 34998 89786
rect 35050 89734 35062 89786
rect 35114 89734 35126 89786
rect 35178 89734 35190 89786
rect 35242 89734 65654 89786
rect 65706 89734 65718 89786
rect 65770 89734 65782 89786
rect 65834 89734 65846 89786
rect 65898 89734 65910 89786
rect 65962 89734 96374 89786
rect 96426 89734 96438 89786
rect 96490 89734 96502 89786
rect 96554 89734 96566 89786
rect 96618 89734 96630 89786
rect 96682 89734 100832 89786
rect 1104 89712 100832 89734
rect 1104 89242 100832 89264
rect 1104 89190 4874 89242
rect 4926 89190 4938 89242
rect 4990 89190 5002 89242
rect 5054 89190 5066 89242
rect 5118 89190 5130 89242
rect 5182 89190 35594 89242
rect 35646 89190 35658 89242
rect 35710 89190 35722 89242
rect 35774 89190 35786 89242
rect 35838 89190 35850 89242
rect 35902 89190 66314 89242
rect 66366 89190 66378 89242
rect 66430 89190 66442 89242
rect 66494 89190 66506 89242
rect 66558 89190 66570 89242
rect 66622 89190 97034 89242
rect 97086 89190 97098 89242
rect 97150 89190 97162 89242
rect 97214 89190 97226 89242
rect 97278 89190 97290 89242
rect 97342 89190 100832 89242
rect 1104 89168 100832 89190
rect 1104 88698 100832 88720
rect 1104 88646 4214 88698
rect 4266 88646 4278 88698
rect 4330 88646 4342 88698
rect 4394 88646 4406 88698
rect 4458 88646 4470 88698
rect 4522 88646 34934 88698
rect 34986 88646 34998 88698
rect 35050 88646 35062 88698
rect 35114 88646 35126 88698
rect 35178 88646 35190 88698
rect 35242 88646 65654 88698
rect 65706 88646 65718 88698
rect 65770 88646 65782 88698
rect 65834 88646 65846 88698
rect 65898 88646 65910 88698
rect 65962 88646 96374 88698
rect 96426 88646 96438 88698
rect 96490 88646 96502 88698
rect 96554 88646 96566 88698
rect 96618 88646 96630 88698
rect 96682 88646 100832 88698
rect 1104 88624 100832 88646
rect 1104 88154 100832 88176
rect 1104 88102 4874 88154
rect 4926 88102 4938 88154
rect 4990 88102 5002 88154
rect 5054 88102 5066 88154
rect 5118 88102 5130 88154
rect 5182 88102 35594 88154
rect 35646 88102 35658 88154
rect 35710 88102 35722 88154
rect 35774 88102 35786 88154
rect 35838 88102 35850 88154
rect 35902 88102 66314 88154
rect 66366 88102 66378 88154
rect 66430 88102 66442 88154
rect 66494 88102 66506 88154
rect 66558 88102 66570 88154
rect 66622 88102 97034 88154
rect 97086 88102 97098 88154
rect 97150 88102 97162 88154
rect 97214 88102 97226 88154
rect 97278 88102 97290 88154
rect 97342 88102 100832 88154
rect 1104 88080 100832 88102
rect 1104 87610 100832 87632
rect 1104 87558 4214 87610
rect 4266 87558 4278 87610
rect 4330 87558 4342 87610
rect 4394 87558 4406 87610
rect 4458 87558 4470 87610
rect 4522 87558 34934 87610
rect 34986 87558 34998 87610
rect 35050 87558 35062 87610
rect 35114 87558 35126 87610
rect 35178 87558 35190 87610
rect 35242 87558 65654 87610
rect 65706 87558 65718 87610
rect 65770 87558 65782 87610
rect 65834 87558 65846 87610
rect 65898 87558 65910 87610
rect 65962 87558 96374 87610
rect 96426 87558 96438 87610
rect 96490 87558 96502 87610
rect 96554 87558 96566 87610
rect 96618 87558 96630 87610
rect 96682 87558 100832 87610
rect 1104 87536 100832 87558
rect 1104 87066 100832 87088
rect 1104 87014 4874 87066
rect 4926 87014 4938 87066
rect 4990 87014 5002 87066
rect 5054 87014 5066 87066
rect 5118 87014 5130 87066
rect 5182 87014 35594 87066
rect 35646 87014 35658 87066
rect 35710 87014 35722 87066
rect 35774 87014 35786 87066
rect 35838 87014 35850 87066
rect 35902 87014 66314 87066
rect 66366 87014 66378 87066
rect 66430 87014 66442 87066
rect 66494 87014 66506 87066
rect 66558 87014 66570 87066
rect 66622 87014 97034 87066
rect 97086 87014 97098 87066
rect 97150 87014 97162 87066
rect 97214 87014 97226 87066
rect 97278 87014 97290 87066
rect 97342 87014 100832 87066
rect 1104 86992 100832 87014
rect 1104 86522 100832 86544
rect 1104 86470 4214 86522
rect 4266 86470 4278 86522
rect 4330 86470 4342 86522
rect 4394 86470 4406 86522
rect 4458 86470 4470 86522
rect 4522 86470 34934 86522
rect 34986 86470 34998 86522
rect 35050 86470 35062 86522
rect 35114 86470 35126 86522
rect 35178 86470 35190 86522
rect 35242 86470 65654 86522
rect 65706 86470 65718 86522
rect 65770 86470 65782 86522
rect 65834 86470 65846 86522
rect 65898 86470 65910 86522
rect 65962 86470 96374 86522
rect 96426 86470 96438 86522
rect 96490 86470 96502 86522
rect 96554 86470 96566 86522
rect 96618 86470 96630 86522
rect 96682 86470 100832 86522
rect 1104 86448 100832 86470
rect 1104 85978 100832 86000
rect 1104 85926 4874 85978
rect 4926 85926 4938 85978
rect 4990 85926 5002 85978
rect 5054 85926 5066 85978
rect 5118 85926 5130 85978
rect 5182 85926 35594 85978
rect 35646 85926 35658 85978
rect 35710 85926 35722 85978
rect 35774 85926 35786 85978
rect 35838 85926 35850 85978
rect 35902 85926 66314 85978
rect 66366 85926 66378 85978
rect 66430 85926 66442 85978
rect 66494 85926 66506 85978
rect 66558 85926 66570 85978
rect 66622 85926 97034 85978
rect 97086 85926 97098 85978
rect 97150 85926 97162 85978
rect 97214 85926 97226 85978
rect 97278 85926 97290 85978
rect 97342 85926 100832 85978
rect 1104 85904 100832 85926
rect 1104 85434 100832 85456
rect 1104 85382 4214 85434
rect 4266 85382 4278 85434
rect 4330 85382 4342 85434
rect 4394 85382 4406 85434
rect 4458 85382 4470 85434
rect 4522 85382 34934 85434
rect 34986 85382 34998 85434
rect 35050 85382 35062 85434
rect 35114 85382 35126 85434
rect 35178 85382 35190 85434
rect 35242 85382 65654 85434
rect 65706 85382 65718 85434
rect 65770 85382 65782 85434
rect 65834 85382 65846 85434
rect 65898 85382 65910 85434
rect 65962 85382 96374 85434
rect 96426 85382 96438 85434
rect 96490 85382 96502 85434
rect 96554 85382 96566 85434
rect 96618 85382 96630 85434
rect 96682 85382 100832 85434
rect 1104 85360 100832 85382
rect 1104 84890 100832 84912
rect 1104 84838 4874 84890
rect 4926 84838 4938 84890
rect 4990 84838 5002 84890
rect 5054 84838 5066 84890
rect 5118 84838 5130 84890
rect 5182 84838 35594 84890
rect 35646 84838 35658 84890
rect 35710 84838 35722 84890
rect 35774 84838 35786 84890
rect 35838 84838 35850 84890
rect 35902 84838 66314 84890
rect 66366 84838 66378 84890
rect 66430 84838 66442 84890
rect 66494 84838 66506 84890
rect 66558 84838 66570 84890
rect 66622 84838 97034 84890
rect 97086 84838 97098 84890
rect 97150 84838 97162 84890
rect 97214 84838 97226 84890
rect 97278 84838 97290 84890
rect 97342 84838 100832 84890
rect 1104 84816 100832 84838
rect 1104 84346 100832 84368
rect 1104 84294 4214 84346
rect 4266 84294 4278 84346
rect 4330 84294 4342 84346
rect 4394 84294 4406 84346
rect 4458 84294 4470 84346
rect 4522 84294 34934 84346
rect 34986 84294 34998 84346
rect 35050 84294 35062 84346
rect 35114 84294 35126 84346
rect 35178 84294 35190 84346
rect 35242 84294 65654 84346
rect 65706 84294 65718 84346
rect 65770 84294 65782 84346
rect 65834 84294 65846 84346
rect 65898 84294 65910 84346
rect 65962 84294 96374 84346
rect 96426 84294 96438 84346
rect 96490 84294 96502 84346
rect 96554 84294 96566 84346
rect 96618 84294 96630 84346
rect 96682 84294 100832 84346
rect 1104 84272 100832 84294
rect 1104 83802 100832 83824
rect 1104 83750 4874 83802
rect 4926 83750 4938 83802
rect 4990 83750 5002 83802
rect 5054 83750 5066 83802
rect 5118 83750 5130 83802
rect 5182 83750 35594 83802
rect 35646 83750 35658 83802
rect 35710 83750 35722 83802
rect 35774 83750 35786 83802
rect 35838 83750 35850 83802
rect 35902 83750 66314 83802
rect 66366 83750 66378 83802
rect 66430 83750 66442 83802
rect 66494 83750 66506 83802
rect 66558 83750 66570 83802
rect 66622 83750 97034 83802
rect 97086 83750 97098 83802
rect 97150 83750 97162 83802
rect 97214 83750 97226 83802
rect 97278 83750 97290 83802
rect 97342 83750 100832 83802
rect 1104 83728 100832 83750
rect 1104 83258 100832 83280
rect 1104 83206 4214 83258
rect 4266 83206 4278 83258
rect 4330 83206 4342 83258
rect 4394 83206 4406 83258
rect 4458 83206 4470 83258
rect 4522 83206 34934 83258
rect 34986 83206 34998 83258
rect 35050 83206 35062 83258
rect 35114 83206 35126 83258
rect 35178 83206 35190 83258
rect 35242 83206 65654 83258
rect 65706 83206 65718 83258
rect 65770 83206 65782 83258
rect 65834 83206 65846 83258
rect 65898 83206 65910 83258
rect 65962 83206 96374 83258
rect 96426 83206 96438 83258
rect 96490 83206 96502 83258
rect 96554 83206 96566 83258
rect 96618 83206 96630 83258
rect 96682 83206 100832 83258
rect 1104 83184 100832 83206
rect 1104 82714 100832 82736
rect 1104 82662 4874 82714
rect 4926 82662 4938 82714
rect 4990 82662 5002 82714
rect 5054 82662 5066 82714
rect 5118 82662 5130 82714
rect 5182 82662 35594 82714
rect 35646 82662 35658 82714
rect 35710 82662 35722 82714
rect 35774 82662 35786 82714
rect 35838 82662 35850 82714
rect 35902 82662 66314 82714
rect 66366 82662 66378 82714
rect 66430 82662 66442 82714
rect 66494 82662 66506 82714
rect 66558 82662 66570 82714
rect 66622 82662 97034 82714
rect 97086 82662 97098 82714
rect 97150 82662 97162 82714
rect 97214 82662 97226 82714
rect 97278 82662 97290 82714
rect 97342 82662 100832 82714
rect 1104 82640 100832 82662
rect 1104 82170 100832 82192
rect 1104 82118 4214 82170
rect 4266 82118 4278 82170
rect 4330 82118 4342 82170
rect 4394 82118 4406 82170
rect 4458 82118 4470 82170
rect 4522 82118 34934 82170
rect 34986 82118 34998 82170
rect 35050 82118 35062 82170
rect 35114 82118 35126 82170
rect 35178 82118 35190 82170
rect 35242 82118 65654 82170
rect 65706 82118 65718 82170
rect 65770 82118 65782 82170
rect 65834 82118 65846 82170
rect 65898 82118 65910 82170
rect 65962 82118 96374 82170
rect 96426 82118 96438 82170
rect 96490 82118 96502 82170
rect 96554 82118 96566 82170
rect 96618 82118 96630 82170
rect 96682 82118 100832 82170
rect 1104 82096 100832 82118
rect 1104 81626 100832 81648
rect 1104 81574 4874 81626
rect 4926 81574 4938 81626
rect 4990 81574 5002 81626
rect 5054 81574 5066 81626
rect 5118 81574 5130 81626
rect 5182 81574 35594 81626
rect 35646 81574 35658 81626
rect 35710 81574 35722 81626
rect 35774 81574 35786 81626
rect 35838 81574 35850 81626
rect 35902 81574 66314 81626
rect 66366 81574 66378 81626
rect 66430 81574 66442 81626
rect 66494 81574 66506 81626
rect 66558 81574 66570 81626
rect 66622 81574 97034 81626
rect 97086 81574 97098 81626
rect 97150 81574 97162 81626
rect 97214 81574 97226 81626
rect 97278 81574 97290 81626
rect 97342 81574 100832 81626
rect 1104 81552 100832 81574
rect 1104 81082 100832 81104
rect 1104 81030 4214 81082
rect 4266 81030 4278 81082
rect 4330 81030 4342 81082
rect 4394 81030 4406 81082
rect 4458 81030 4470 81082
rect 4522 81030 34934 81082
rect 34986 81030 34998 81082
rect 35050 81030 35062 81082
rect 35114 81030 35126 81082
rect 35178 81030 35190 81082
rect 35242 81030 65654 81082
rect 65706 81030 65718 81082
rect 65770 81030 65782 81082
rect 65834 81030 65846 81082
rect 65898 81030 65910 81082
rect 65962 81030 96374 81082
rect 96426 81030 96438 81082
rect 96490 81030 96502 81082
rect 96554 81030 96566 81082
rect 96618 81030 96630 81082
rect 96682 81030 100832 81082
rect 1104 81008 100832 81030
rect 1104 80538 100832 80560
rect 1104 80486 4874 80538
rect 4926 80486 4938 80538
rect 4990 80486 5002 80538
rect 5054 80486 5066 80538
rect 5118 80486 5130 80538
rect 5182 80486 35594 80538
rect 35646 80486 35658 80538
rect 35710 80486 35722 80538
rect 35774 80486 35786 80538
rect 35838 80486 35850 80538
rect 35902 80486 66314 80538
rect 66366 80486 66378 80538
rect 66430 80486 66442 80538
rect 66494 80486 66506 80538
rect 66558 80486 66570 80538
rect 66622 80486 97034 80538
rect 97086 80486 97098 80538
rect 97150 80486 97162 80538
rect 97214 80486 97226 80538
rect 97278 80486 97290 80538
rect 97342 80486 100832 80538
rect 1104 80464 100832 80486
rect 1104 79994 100832 80016
rect 1104 79942 4214 79994
rect 4266 79942 4278 79994
rect 4330 79942 4342 79994
rect 4394 79942 4406 79994
rect 4458 79942 4470 79994
rect 4522 79942 34934 79994
rect 34986 79942 34998 79994
rect 35050 79942 35062 79994
rect 35114 79942 35126 79994
rect 35178 79942 35190 79994
rect 35242 79942 65654 79994
rect 65706 79942 65718 79994
rect 65770 79942 65782 79994
rect 65834 79942 65846 79994
rect 65898 79942 65910 79994
rect 65962 79942 96374 79994
rect 96426 79942 96438 79994
rect 96490 79942 96502 79994
rect 96554 79942 96566 79994
rect 96618 79942 96630 79994
rect 96682 79942 100832 79994
rect 1104 79920 100832 79942
rect 1104 79450 100832 79472
rect 1104 79398 4874 79450
rect 4926 79398 4938 79450
rect 4990 79398 5002 79450
rect 5054 79398 5066 79450
rect 5118 79398 5130 79450
rect 5182 79398 35594 79450
rect 35646 79398 35658 79450
rect 35710 79398 35722 79450
rect 35774 79398 35786 79450
rect 35838 79398 35850 79450
rect 35902 79398 66314 79450
rect 66366 79398 66378 79450
rect 66430 79398 66442 79450
rect 66494 79398 66506 79450
rect 66558 79398 66570 79450
rect 66622 79398 97034 79450
rect 97086 79398 97098 79450
rect 97150 79398 97162 79450
rect 97214 79398 97226 79450
rect 97278 79398 97290 79450
rect 97342 79398 100832 79450
rect 1104 79376 100832 79398
rect 1104 78906 100832 78928
rect 1104 78854 4214 78906
rect 4266 78854 4278 78906
rect 4330 78854 4342 78906
rect 4394 78854 4406 78906
rect 4458 78854 4470 78906
rect 4522 78854 34934 78906
rect 34986 78854 34998 78906
rect 35050 78854 35062 78906
rect 35114 78854 35126 78906
rect 35178 78854 35190 78906
rect 35242 78854 65654 78906
rect 65706 78854 65718 78906
rect 65770 78854 65782 78906
rect 65834 78854 65846 78906
rect 65898 78854 65910 78906
rect 65962 78854 96374 78906
rect 96426 78854 96438 78906
rect 96490 78854 96502 78906
rect 96554 78854 96566 78906
rect 96618 78854 96630 78906
rect 96682 78854 100832 78906
rect 1104 78832 100832 78854
rect 1104 78362 100832 78384
rect 1104 78310 4874 78362
rect 4926 78310 4938 78362
rect 4990 78310 5002 78362
rect 5054 78310 5066 78362
rect 5118 78310 5130 78362
rect 5182 78310 35594 78362
rect 35646 78310 35658 78362
rect 35710 78310 35722 78362
rect 35774 78310 35786 78362
rect 35838 78310 35850 78362
rect 35902 78310 66314 78362
rect 66366 78310 66378 78362
rect 66430 78310 66442 78362
rect 66494 78310 66506 78362
rect 66558 78310 66570 78362
rect 66622 78310 97034 78362
rect 97086 78310 97098 78362
rect 97150 78310 97162 78362
rect 97214 78310 97226 78362
rect 97278 78310 97290 78362
rect 97342 78310 100832 78362
rect 1104 78288 100832 78310
rect 1104 77818 100832 77840
rect 1104 77766 4214 77818
rect 4266 77766 4278 77818
rect 4330 77766 4342 77818
rect 4394 77766 4406 77818
rect 4458 77766 4470 77818
rect 4522 77766 34934 77818
rect 34986 77766 34998 77818
rect 35050 77766 35062 77818
rect 35114 77766 35126 77818
rect 35178 77766 35190 77818
rect 35242 77766 65654 77818
rect 65706 77766 65718 77818
rect 65770 77766 65782 77818
rect 65834 77766 65846 77818
rect 65898 77766 65910 77818
rect 65962 77766 96374 77818
rect 96426 77766 96438 77818
rect 96490 77766 96502 77818
rect 96554 77766 96566 77818
rect 96618 77766 96630 77818
rect 96682 77766 100832 77818
rect 1104 77744 100832 77766
rect 43530 77664 43536 77716
rect 43588 77664 43594 77716
rect 47486 77664 47492 77716
rect 47544 77664 47550 77716
rect 49694 77664 49700 77716
rect 49752 77664 49758 77716
rect 53098 77664 53104 77716
rect 53156 77664 53162 77716
rect 55122 77664 55128 77716
rect 55180 77664 55186 77716
rect 57330 77664 57336 77716
rect 57388 77664 57394 77716
rect 59170 77664 59176 77716
rect 59228 77664 59234 77716
rect 41785 77571 41843 77577
rect 41785 77537 41797 77571
rect 41831 77568 41843 77571
rect 43622 77568 43628 77580
rect 41831 77540 43628 77568
rect 41831 77537 41843 77540
rect 41785 77531 41843 77537
rect 43622 77528 43628 77540
rect 43680 77568 43686 77580
rect 45741 77571 45799 77577
rect 45741 77568 45753 77571
rect 43680 77540 45753 77568
rect 43680 77528 43686 77540
rect 45741 77537 45753 77540
rect 45787 77568 45799 77571
rect 47949 77571 48007 77577
rect 47949 77568 47961 77571
rect 45787 77540 47961 77568
rect 45787 77537 45799 77540
rect 45741 77531 45799 77537
rect 47949 77537 47961 77540
rect 47995 77568 48007 77571
rect 49418 77568 49424 77580
rect 47995 77540 49424 77568
rect 47995 77537 48007 77540
rect 47949 77531 48007 77537
rect 49418 77528 49424 77540
rect 49476 77568 49482 77580
rect 51353 77571 51411 77577
rect 51353 77568 51365 77571
rect 49476 77540 51365 77568
rect 49476 77528 49482 77540
rect 51353 77537 51365 77540
rect 51399 77568 51411 77571
rect 53377 77571 53435 77577
rect 53377 77568 53389 77571
rect 51399 77540 53389 77568
rect 51399 77537 51411 77540
rect 51353 77531 51411 77537
rect 53377 77537 53389 77540
rect 53423 77568 53435 77571
rect 55585 77571 55643 77577
rect 55585 77568 55597 77571
rect 53423 77540 55597 77568
rect 53423 77537 53435 77540
rect 53377 77531 53435 77537
rect 55585 77537 55597 77540
rect 55631 77568 55643 77571
rect 57425 77571 57483 77577
rect 57425 77568 57437 77571
rect 55631 77540 57437 77568
rect 55631 77537 55643 77540
rect 55585 77531 55643 77537
rect 57425 77537 57437 77540
rect 57471 77537 57483 77571
rect 57425 77531 57483 77537
rect 42061 77435 42119 77441
rect 42061 77401 42073 77435
rect 42107 77401 42119 77435
rect 45646 77432 45652 77444
rect 43286 77404 45652 77432
rect 42061 77395 42119 77401
rect 41693 77367 41751 77373
rect 41693 77333 41705 77367
rect 41739 77364 41751 77367
rect 41782 77364 41788 77376
rect 41739 77336 41788 77364
rect 41739 77333 41751 77336
rect 41693 77327 41751 77333
rect 41782 77324 41788 77336
rect 41840 77364 41846 77376
rect 42076 77364 42104 77395
rect 45646 77392 45652 77404
rect 45704 77392 45710 77444
rect 45738 77392 45744 77444
rect 45796 77432 45802 77444
rect 46017 77435 46075 77441
rect 46017 77432 46029 77435
rect 45796 77404 46029 77432
rect 45796 77392 45802 77404
rect 46017 77401 46029 77404
rect 46063 77401 46075 77435
rect 47242 77404 47900 77432
rect 46017 77395 46075 77401
rect 41840 77336 42104 77364
rect 47872 77364 47900 77404
rect 47946 77392 47952 77444
rect 48004 77432 48010 77444
rect 48225 77435 48283 77441
rect 48225 77432 48237 77435
rect 48004 77404 48237 77432
rect 48004 77392 48010 77404
rect 48225 77401 48237 77404
rect 48271 77401 48283 77435
rect 51074 77432 51080 77444
rect 49450 77404 51080 77432
rect 48225 77395 48283 77401
rect 51074 77392 51080 77404
rect 51132 77392 51138 77444
rect 51258 77392 51264 77444
rect 51316 77432 51322 77444
rect 51629 77435 51687 77441
rect 51629 77432 51641 77435
rect 51316 77404 51641 77432
rect 51316 77392 51322 77404
rect 51629 77401 51641 77404
rect 51675 77401 51687 77435
rect 53374 77432 53380 77444
rect 52854 77404 53380 77432
rect 51629 77395 51687 77401
rect 53374 77392 53380 77404
rect 53432 77392 53438 77444
rect 53653 77435 53711 77441
rect 53653 77401 53665 77435
rect 53699 77401 53711 77435
rect 54878 77404 55214 77432
rect 53653 77395 53711 77401
rect 49970 77364 49976 77376
rect 47872 77336 49976 77364
rect 41840 77324 41846 77336
rect 49970 77324 49976 77336
rect 50028 77324 50034 77376
rect 53282 77324 53288 77376
rect 53340 77364 53346 77376
rect 53668 77364 53696 77395
rect 53340 77336 53696 77364
rect 55186 77364 55214 77404
rect 55582 77392 55588 77444
rect 55640 77432 55646 77444
rect 55861 77435 55919 77441
rect 55861 77432 55873 77435
rect 55640 77404 55873 77432
rect 55640 77392 55646 77404
rect 55861 77401 55873 77404
rect 55907 77401 55919 77435
rect 57422 77432 57428 77444
rect 57086 77404 57428 77432
rect 55861 77395 55919 77401
rect 57422 77392 57428 77404
rect 57480 77392 57486 77444
rect 57701 77435 57759 77441
rect 57701 77432 57713 77435
rect 57532 77404 57713 77432
rect 57532 77376 57560 77404
rect 57701 77401 57713 77404
rect 57747 77401 57759 77435
rect 59262 77432 59268 77444
rect 58926 77404 59268 77432
rect 57701 77395 57759 77401
rect 59262 77392 59268 77404
rect 59320 77392 59326 77444
rect 56870 77364 56876 77376
rect 55186 77336 56876 77364
rect 53340 77324 53346 77336
rect 56870 77324 56876 77336
rect 56928 77324 56934 77376
rect 57514 77324 57520 77376
rect 57572 77324 57578 77376
rect 1104 77274 100832 77296
rect 1104 77222 4874 77274
rect 4926 77222 4938 77274
rect 4990 77222 5002 77274
rect 5054 77222 5066 77274
rect 5118 77222 5130 77274
rect 5182 77222 35594 77274
rect 35646 77222 35658 77274
rect 35710 77222 35722 77274
rect 35774 77222 35786 77274
rect 35838 77222 35850 77274
rect 35902 77222 66314 77274
rect 66366 77222 66378 77274
rect 66430 77222 66442 77274
rect 66494 77222 66506 77274
rect 66558 77222 66570 77274
rect 66622 77222 97034 77274
rect 97086 77222 97098 77274
rect 97150 77222 97162 77274
rect 97214 77222 97226 77274
rect 97278 77222 97290 77274
rect 97342 77222 100832 77274
rect 1104 77200 100832 77222
rect 45370 77120 45376 77172
rect 45428 77120 45434 77172
rect 51166 77120 51172 77172
rect 51224 77120 51230 77172
rect 48222 77092 48228 77104
rect 45126 77064 48228 77092
rect 48222 77052 48228 77064
rect 48280 77052 48286 77104
rect 49602 77052 49608 77104
rect 49660 77092 49666 77104
rect 49697 77095 49755 77101
rect 49697 77092 49709 77095
rect 49660 77064 49709 77092
rect 49660 77052 49666 77064
rect 49697 77061 49709 77064
rect 49743 77061 49755 77095
rect 53190 77092 53196 77104
rect 50922 77064 53196 77092
rect 49697 77055 49755 77061
rect 53190 77052 53196 77064
rect 53248 77052 53254 77104
rect 43622 76984 43628 77036
rect 43680 76984 43686 77036
rect 49418 76984 49424 77036
rect 49476 76984 49482 77036
rect 43901 76959 43959 76965
rect 43901 76956 43913 76959
rect 43640 76928 43913 76956
rect 43640 76900 43668 76928
rect 43901 76925 43913 76928
rect 43947 76925 43959 76959
rect 43901 76919 43959 76925
rect 43622 76848 43628 76900
rect 43680 76848 43686 76900
rect 41782 76780 41788 76832
rect 41840 76780 41846 76832
rect 45738 76780 45744 76832
rect 45796 76780 45802 76832
rect 47946 76780 47952 76832
rect 48004 76780 48010 76832
rect 51258 76780 51264 76832
rect 51316 76820 51322 76832
rect 51353 76823 51411 76829
rect 51353 76820 51365 76823
rect 51316 76792 51365 76820
rect 51316 76780 51322 76792
rect 51353 76789 51365 76792
rect 51399 76789 51411 76823
rect 51353 76783 51411 76789
rect 53282 76780 53288 76832
rect 53340 76820 53346 76832
rect 53377 76823 53435 76829
rect 53377 76820 53389 76823
rect 53340 76792 53389 76820
rect 53340 76780 53346 76792
rect 53377 76789 53389 76792
rect 53423 76789 53435 76823
rect 53377 76783 53435 76789
rect 55582 76780 55588 76832
rect 55640 76780 55646 76832
rect 57514 76780 57520 76832
rect 57572 76780 57578 76832
rect 1104 76730 100832 76752
rect 1104 76678 4214 76730
rect 4266 76678 4278 76730
rect 4330 76678 4342 76730
rect 4394 76678 4406 76730
rect 4458 76678 4470 76730
rect 4522 76678 34934 76730
rect 34986 76678 34998 76730
rect 35050 76678 35062 76730
rect 35114 76678 35126 76730
rect 35178 76678 35190 76730
rect 35242 76678 65654 76730
rect 65706 76678 65718 76730
rect 65770 76678 65782 76730
rect 65834 76678 65846 76730
rect 65898 76678 65910 76730
rect 65962 76678 96374 76730
rect 96426 76678 96438 76730
rect 96490 76678 96502 76730
rect 96554 76678 96566 76730
rect 96618 76678 96630 76730
rect 96682 76678 100832 76730
rect 1104 76656 100832 76678
rect 49513 76619 49571 76625
rect 49513 76585 49525 76619
rect 49559 76616 49571 76619
rect 49602 76616 49608 76628
rect 49559 76588 49608 76616
rect 49559 76585 49571 76588
rect 49513 76579 49571 76585
rect 49602 76576 49608 76588
rect 49660 76576 49666 76628
rect 43622 76236 43628 76288
rect 43680 76236 43686 76288
rect 1104 76186 100832 76208
rect 1104 76134 4874 76186
rect 4926 76134 4938 76186
rect 4990 76134 5002 76186
rect 5054 76134 5066 76186
rect 5118 76134 5130 76186
rect 5182 76134 35594 76186
rect 35646 76134 35658 76186
rect 35710 76134 35722 76186
rect 35774 76134 35786 76186
rect 35838 76134 35850 76186
rect 35902 76134 66314 76186
rect 66366 76134 66378 76186
rect 66430 76134 66442 76186
rect 66494 76134 66506 76186
rect 66558 76134 66570 76186
rect 66622 76134 97034 76186
rect 97086 76134 97098 76186
rect 97150 76134 97162 76186
rect 97214 76134 97226 76186
rect 97278 76134 97290 76186
rect 97342 76134 100832 76186
rect 1104 76112 100832 76134
rect 1104 75642 100832 75664
rect 1104 75590 4214 75642
rect 4266 75590 4278 75642
rect 4330 75590 4342 75642
rect 4394 75590 4406 75642
rect 4458 75590 4470 75642
rect 4522 75590 34934 75642
rect 34986 75590 34998 75642
rect 35050 75590 35062 75642
rect 35114 75590 35126 75642
rect 35178 75590 35190 75642
rect 35242 75590 65654 75642
rect 65706 75590 65718 75642
rect 65770 75590 65782 75642
rect 65834 75590 65846 75642
rect 65898 75590 65910 75642
rect 65962 75590 96374 75642
rect 96426 75590 96438 75642
rect 96490 75590 96502 75642
rect 96554 75590 96566 75642
rect 96618 75590 96630 75642
rect 96682 75590 100832 75642
rect 1104 75568 100832 75590
rect 1104 75098 100832 75120
rect 1104 75046 4874 75098
rect 4926 75046 4938 75098
rect 4990 75046 5002 75098
rect 5054 75046 5066 75098
rect 5118 75046 5130 75098
rect 5182 75046 35594 75098
rect 35646 75046 35658 75098
rect 35710 75046 35722 75098
rect 35774 75046 35786 75098
rect 35838 75046 35850 75098
rect 35902 75046 66314 75098
rect 66366 75046 66378 75098
rect 66430 75046 66442 75098
rect 66494 75046 66506 75098
rect 66558 75046 66570 75098
rect 66622 75046 97034 75098
rect 97086 75046 97098 75098
rect 97150 75046 97162 75098
rect 97214 75046 97226 75098
rect 97278 75046 97290 75098
rect 97342 75046 100832 75098
rect 1104 75024 100832 75046
rect 45646 74944 45652 74996
rect 45704 74984 45710 74996
rect 46569 74987 46627 74993
rect 46569 74984 46581 74987
rect 45704 74956 46581 74984
rect 45704 74944 45710 74956
rect 46569 74953 46581 74956
rect 46615 74953 46627 74987
rect 46569 74947 46627 74953
rect 48222 74944 48228 74996
rect 48280 74944 48286 74996
rect 49970 74944 49976 74996
rect 50028 74944 50034 74996
rect 51074 74944 51080 74996
rect 51132 74984 51138 74996
rect 51905 74987 51963 74993
rect 51905 74984 51917 74987
rect 51132 74956 51917 74984
rect 51132 74944 51138 74956
rect 51905 74953 51917 74956
rect 51951 74953 51963 74987
rect 51905 74947 51963 74953
rect 53190 74944 53196 74996
rect 53248 74944 53254 74996
rect 53374 74944 53380 74996
rect 53432 74984 53438 74996
rect 54849 74987 54907 74993
rect 54849 74984 54861 74987
rect 53432 74956 54861 74984
rect 53432 74944 53438 74956
rect 54849 74953 54861 74956
rect 54895 74953 54907 74987
rect 54849 74947 54907 74953
rect 56870 74944 56876 74996
rect 56928 74944 56934 74996
rect 57422 74944 57428 74996
rect 57480 74984 57486 74996
rect 58345 74987 58403 74993
rect 58345 74984 58357 74987
rect 57480 74956 58357 74984
rect 57480 74944 57486 74956
rect 58345 74953 58357 74956
rect 58391 74953 58403 74987
rect 58345 74947 58403 74953
rect 59262 74944 59268 74996
rect 59320 74984 59326 74996
rect 60645 74987 60703 74993
rect 60645 74984 60657 74987
rect 59320 74956 60657 74984
rect 59320 74944 59326 74956
rect 60645 74953 60657 74956
rect 60691 74953 60703 74987
rect 60645 74947 60703 74953
rect 50080 74888 53328 74916
rect 46658 74808 46664 74860
rect 46716 74848 46722 74860
rect 50080 74857 50108 74888
rect 53300 74857 53328 74888
rect 60200 74888 60596 74916
rect 60200 74857 60228 74888
rect 60568 74857 60596 74888
rect 48317 74851 48375 74857
rect 48317 74848 48329 74851
rect 46716 74820 48329 74848
rect 46716 74808 46722 74820
rect 48317 74817 48329 74820
rect 48363 74848 48375 74851
rect 50065 74851 50123 74857
rect 50065 74848 50077 74851
rect 48363 74820 50077 74848
rect 48363 74817 48375 74820
rect 48317 74811 48375 74817
rect 50065 74817 50077 74820
rect 50111 74817 50123 74851
rect 50065 74811 50123 74817
rect 51997 74851 52055 74857
rect 51997 74817 52009 74851
rect 52043 74817 52055 74851
rect 51997 74811 52055 74817
rect 53285 74851 53343 74857
rect 53285 74817 53297 74851
rect 53331 74848 53343 74851
rect 54941 74851 54999 74857
rect 54941 74848 54953 74851
rect 53331 74820 54953 74848
rect 53331 74817 53343 74820
rect 53285 74811 53343 74817
rect 54941 74817 54953 74820
rect 54987 74848 54999 74851
rect 56965 74851 57023 74857
rect 56965 74848 56977 74851
rect 54987 74820 56977 74848
rect 54987 74817 54999 74820
rect 54941 74811 54999 74817
rect 56965 74817 56977 74820
rect 57011 74848 57023 74851
rect 58437 74851 58495 74857
rect 58437 74848 58449 74851
rect 57011 74820 58449 74848
rect 57011 74817 57023 74820
rect 56965 74811 57023 74817
rect 58437 74817 58449 74820
rect 58483 74848 58495 74851
rect 60185 74851 60243 74857
rect 60185 74848 60197 74851
rect 58483 74820 60197 74848
rect 58483 74817 58495 74820
rect 58437 74811 58495 74817
rect 60185 74817 60197 74820
rect 60231 74817 60243 74851
rect 60185 74811 60243 74817
rect 60461 74851 60519 74857
rect 60461 74817 60473 74851
rect 60507 74817 60519 74851
rect 60461 74811 60519 74817
rect 60553 74851 60611 74857
rect 60553 74817 60565 74851
rect 60599 74817 60611 74851
rect 83918 74848 83924 74860
rect 60553 74811 60611 74817
rect 64846 74820 83924 74848
rect 52012 74780 52040 74811
rect 60476 74780 60504 74811
rect 64846 74780 64874 74820
rect 83918 74808 83924 74820
rect 83976 74808 83982 74860
rect 52012 74752 64874 74780
rect 1104 74554 100832 74576
rect 1104 74502 4214 74554
rect 4266 74502 4278 74554
rect 4330 74502 4342 74554
rect 4394 74502 4406 74554
rect 4458 74502 4470 74554
rect 4522 74502 34934 74554
rect 34986 74502 34998 74554
rect 35050 74502 35062 74554
rect 35114 74502 35126 74554
rect 35178 74502 35190 74554
rect 35242 74502 65654 74554
rect 65706 74502 65718 74554
rect 65770 74502 65782 74554
rect 65834 74502 65846 74554
rect 65898 74502 65910 74554
rect 65962 74502 96374 74554
rect 96426 74502 96438 74554
rect 96490 74502 96502 74554
rect 96554 74502 96566 74554
rect 96618 74502 96630 74554
rect 96682 74502 100832 74554
rect 1104 74480 100832 74502
rect 1104 74010 100832 74032
rect 1104 73958 4874 74010
rect 4926 73958 4938 74010
rect 4990 73958 5002 74010
rect 5054 73958 5066 74010
rect 5118 73958 5130 74010
rect 5182 73958 35594 74010
rect 35646 73958 35658 74010
rect 35710 73958 35722 74010
rect 35774 73958 35786 74010
rect 35838 73958 35850 74010
rect 35902 73958 66314 74010
rect 66366 73958 66378 74010
rect 66430 73958 66442 74010
rect 66494 73958 66506 74010
rect 66558 73958 66570 74010
rect 66622 73958 97034 74010
rect 97086 73958 97098 74010
rect 97150 73958 97162 74010
rect 97214 73958 97226 74010
rect 97278 73958 97290 74010
rect 97342 73958 100832 74010
rect 1104 73936 100832 73958
rect 1104 73466 100832 73488
rect 1104 73414 4214 73466
rect 4266 73414 4278 73466
rect 4330 73414 4342 73466
rect 4394 73414 4406 73466
rect 4458 73414 4470 73466
rect 4522 73414 34934 73466
rect 34986 73414 34998 73466
rect 35050 73414 35062 73466
rect 35114 73414 35126 73466
rect 35178 73414 35190 73466
rect 35242 73414 65654 73466
rect 65706 73414 65718 73466
rect 65770 73414 65782 73466
rect 65834 73414 65846 73466
rect 65898 73414 65910 73466
rect 65962 73414 96374 73466
rect 96426 73414 96438 73466
rect 96490 73414 96502 73466
rect 96554 73414 96566 73466
rect 96618 73414 96630 73466
rect 96682 73414 100832 73466
rect 1104 73392 100832 73414
rect 1104 72922 100832 72944
rect 1104 72870 4874 72922
rect 4926 72870 4938 72922
rect 4990 72870 5002 72922
rect 5054 72870 5066 72922
rect 5118 72870 5130 72922
rect 5182 72870 35594 72922
rect 35646 72870 35658 72922
rect 35710 72870 35722 72922
rect 35774 72870 35786 72922
rect 35838 72870 35850 72922
rect 35902 72870 66314 72922
rect 66366 72870 66378 72922
rect 66430 72870 66442 72922
rect 66494 72870 66506 72922
rect 66558 72870 66570 72922
rect 66622 72870 97034 72922
rect 97086 72870 97098 72922
rect 97150 72870 97162 72922
rect 97214 72870 97226 72922
rect 97278 72870 97290 72922
rect 97342 72870 100832 72922
rect 1104 72848 100832 72870
rect 1104 72378 100832 72400
rect 1104 72326 4214 72378
rect 4266 72326 4278 72378
rect 4330 72326 4342 72378
rect 4394 72326 4406 72378
rect 4458 72326 4470 72378
rect 4522 72326 34934 72378
rect 34986 72326 34998 72378
rect 35050 72326 35062 72378
rect 35114 72326 35126 72378
rect 35178 72326 35190 72378
rect 35242 72326 65654 72378
rect 65706 72326 65718 72378
rect 65770 72326 65782 72378
rect 65834 72326 65846 72378
rect 65898 72326 65910 72378
rect 65962 72326 96374 72378
rect 96426 72326 96438 72378
rect 96490 72326 96502 72378
rect 96554 72326 96566 72378
rect 96618 72326 96630 72378
rect 96682 72326 100832 72378
rect 1104 72304 100832 72326
rect 1104 71834 100832 71856
rect 1104 71782 4874 71834
rect 4926 71782 4938 71834
rect 4990 71782 5002 71834
rect 5054 71782 5066 71834
rect 5118 71782 5130 71834
rect 5182 71782 35594 71834
rect 35646 71782 35658 71834
rect 35710 71782 35722 71834
rect 35774 71782 35786 71834
rect 35838 71782 35850 71834
rect 35902 71782 66314 71834
rect 66366 71782 66378 71834
rect 66430 71782 66442 71834
rect 66494 71782 66506 71834
rect 66558 71782 66570 71834
rect 66622 71782 97034 71834
rect 97086 71782 97098 71834
rect 97150 71782 97162 71834
rect 97214 71782 97226 71834
rect 97278 71782 97290 71834
rect 97342 71782 100832 71834
rect 1104 71760 100832 71782
rect 1104 71290 100832 71312
rect 1104 71238 4214 71290
rect 4266 71238 4278 71290
rect 4330 71238 4342 71290
rect 4394 71238 4406 71290
rect 4458 71238 4470 71290
rect 4522 71238 34934 71290
rect 34986 71238 34998 71290
rect 35050 71238 35062 71290
rect 35114 71238 35126 71290
rect 35178 71238 35190 71290
rect 35242 71238 65654 71290
rect 65706 71238 65718 71290
rect 65770 71238 65782 71290
rect 65834 71238 65846 71290
rect 65898 71238 65910 71290
rect 65962 71238 96374 71290
rect 96426 71238 96438 71290
rect 96490 71238 96502 71290
rect 96554 71238 96566 71290
rect 96618 71238 96630 71290
rect 96682 71238 100832 71290
rect 1104 71216 100832 71238
rect 1104 70746 100832 70768
rect 1104 70694 4874 70746
rect 4926 70694 4938 70746
rect 4990 70694 5002 70746
rect 5054 70694 5066 70746
rect 5118 70694 5130 70746
rect 5182 70694 35594 70746
rect 35646 70694 35658 70746
rect 35710 70694 35722 70746
rect 35774 70694 35786 70746
rect 35838 70694 35850 70746
rect 35902 70694 66314 70746
rect 66366 70694 66378 70746
rect 66430 70694 66442 70746
rect 66494 70694 66506 70746
rect 66558 70694 66570 70746
rect 66622 70694 97034 70746
rect 97086 70694 97098 70746
rect 97150 70694 97162 70746
rect 97214 70694 97226 70746
rect 97278 70694 97290 70746
rect 97342 70694 100832 70746
rect 1104 70672 100832 70694
rect 1104 70202 100832 70224
rect 1104 70150 4214 70202
rect 4266 70150 4278 70202
rect 4330 70150 4342 70202
rect 4394 70150 4406 70202
rect 4458 70150 4470 70202
rect 4522 70150 34934 70202
rect 34986 70150 34998 70202
rect 35050 70150 35062 70202
rect 35114 70150 35126 70202
rect 35178 70150 35190 70202
rect 35242 70150 65654 70202
rect 65706 70150 65718 70202
rect 65770 70150 65782 70202
rect 65834 70150 65846 70202
rect 65898 70150 65910 70202
rect 65962 70150 96374 70202
rect 96426 70150 96438 70202
rect 96490 70150 96502 70202
rect 96554 70150 96566 70202
rect 96618 70150 96630 70202
rect 96682 70150 100832 70202
rect 1104 70128 100832 70150
rect 1104 69658 100832 69680
rect 1104 69606 4874 69658
rect 4926 69606 4938 69658
rect 4990 69606 5002 69658
rect 5054 69606 5066 69658
rect 5118 69606 5130 69658
rect 5182 69606 35594 69658
rect 35646 69606 35658 69658
rect 35710 69606 35722 69658
rect 35774 69606 35786 69658
rect 35838 69606 35850 69658
rect 35902 69606 66314 69658
rect 66366 69606 66378 69658
rect 66430 69606 66442 69658
rect 66494 69606 66506 69658
rect 66558 69606 66570 69658
rect 66622 69606 97034 69658
rect 97086 69606 97098 69658
rect 97150 69606 97162 69658
rect 97214 69606 97226 69658
rect 97278 69606 97290 69658
rect 97342 69606 100832 69658
rect 1104 69584 100832 69606
rect 1104 69114 100832 69136
rect 1104 69062 4214 69114
rect 4266 69062 4278 69114
rect 4330 69062 4342 69114
rect 4394 69062 4406 69114
rect 4458 69062 4470 69114
rect 4522 69062 34934 69114
rect 34986 69062 34998 69114
rect 35050 69062 35062 69114
rect 35114 69062 35126 69114
rect 35178 69062 35190 69114
rect 35242 69062 65654 69114
rect 65706 69062 65718 69114
rect 65770 69062 65782 69114
rect 65834 69062 65846 69114
rect 65898 69062 65910 69114
rect 65962 69062 96374 69114
rect 96426 69062 96438 69114
rect 96490 69062 96502 69114
rect 96554 69062 96566 69114
rect 96618 69062 96630 69114
rect 96682 69062 100832 69114
rect 1104 69040 100832 69062
rect 1104 68570 100832 68592
rect 1104 68518 4874 68570
rect 4926 68518 4938 68570
rect 4990 68518 5002 68570
rect 5054 68518 5066 68570
rect 5118 68518 5130 68570
rect 5182 68518 35594 68570
rect 35646 68518 35658 68570
rect 35710 68518 35722 68570
rect 35774 68518 35786 68570
rect 35838 68518 35850 68570
rect 35902 68518 66314 68570
rect 66366 68518 66378 68570
rect 66430 68518 66442 68570
rect 66494 68518 66506 68570
rect 66558 68518 66570 68570
rect 66622 68518 97034 68570
rect 97086 68518 97098 68570
rect 97150 68518 97162 68570
rect 97214 68518 97226 68570
rect 97278 68518 97290 68570
rect 97342 68518 100832 68570
rect 1104 68496 100832 68518
rect 1104 68026 100832 68048
rect 1104 67974 4214 68026
rect 4266 67974 4278 68026
rect 4330 67974 4342 68026
rect 4394 67974 4406 68026
rect 4458 67974 4470 68026
rect 4522 67974 34934 68026
rect 34986 67974 34998 68026
rect 35050 67974 35062 68026
rect 35114 67974 35126 68026
rect 35178 67974 35190 68026
rect 35242 67974 65654 68026
rect 65706 67974 65718 68026
rect 65770 67974 65782 68026
rect 65834 67974 65846 68026
rect 65898 67974 65910 68026
rect 65962 67974 96374 68026
rect 96426 67974 96438 68026
rect 96490 67974 96502 68026
rect 96554 67974 96566 68026
rect 96618 67974 96630 68026
rect 96682 67974 100832 68026
rect 1104 67952 100832 67974
rect 1104 67482 100832 67504
rect 1104 67430 4874 67482
rect 4926 67430 4938 67482
rect 4990 67430 5002 67482
rect 5054 67430 5066 67482
rect 5118 67430 5130 67482
rect 5182 67430 35594 67482
rect 35646 67430 35658 67482
rect 35710 67430 35722 67482
rect 35774 67430 35786 67482
rect 35838 67430 35850 67482
rect 35902 67430 66314 67482
rect 66366 67430 66378 67482
rect 66430 67430 66442 67482
rect 66494 67430 66506 67482
rect 66558 67430 66570 67482
rect 66622 67430 97034 67482
rect 97086 67430 97098 67482
rect 97150 67430 97162 67482
rect 97214 67430 97226 67482
rect 97278 67430 97290 67482
rect 97342 67430 100832 67482
rect 1104 67408 100832 67430
rect 1104 66938 100832 66960
rect 1104 66886 4214 66938
rect 4266 66886 4278 66938
rect 4330 66886 4342 66938
rect 4394 66886 4406 66938
rect 4458 66886 4470 66938
rect 4522 66886 34934 66938
rect 34986 66886 34998 66938
rect 35050 66886 35062 66938
rect 35114 66886 35126 66938
rect 35178 66886 35190 66938
rect 35242 66886 65654 66938
rect 65706 66886 65718 66938
rect 65770 66886 65782 66938
rect 65834 66886 65846 66938
rect 65898 66886 65910 66938
rect 65962 66886 96374 66938
rect 96426 66886 96438 66938
rect 96490 66886 96502 66938
rect 96554 66886 96566 66938
rect 96618 66886 96630 66938
rect 96682 66886 100832 66938
rect 1104 66864 100832 66886
rect 1104 66394 100832 66416
rect 1104 66342 4874 66394
rect 4926 66342 4938 66394
rect 4990 66342 5002 66394
rect 5054 66342 5066 66394
rect 5118 66342 5130 66394
rect 5182 66342 35594 66394
rect 35646 66342 35658 66394
rect 35710 66342 35722 66394
rect 35774 66342 35786 66394
rect 35838 66342 35850 66394
rect 35902 66342 66314 66394
rect 66366 66342 66378 66394
rect 66430 66342 66442 66394
rect 66494 66342 66506 66394
rect 66558 66342 66570 66394
rect 66622 66342 97034 66394
rect 97086 66342 97098 66394
rect 97150 66342 97162 66394
rect 97214 66342 97226 66394
rect 97278 66342 97290 66394
rect 97342 66342 100832 66394
rect 1104 66320 100832 66342
rect 1104 65850 100832 65872
rect 1104 65798 4214 65850
rect 4266 65798 4278 65850
rect 4330 65798 4342 65850
rect 4394 65798 4406 65850
rect 4458 65798 4470 65850
rect 4522 65798 34934 65850
rect 34986 65798 34998 65850
rect 35050 65798 35062 65850
rect 35114 65798 35126 65850
rect 35178 65798 35190 65850
rect 35242 65798 65654 65850
rect 65706 65798 65718 65850
rect 65770 65798 65782 65850
rect 65834 65798 65846 65850
rect 65898 65798 65910 65850
rect 65962 65798 96374 65850
rect 96426 65798 96438 65850
rect 96490 65798 96502 65850
rect 96554 65798 96566 65850
rect 96618 65798 96630 65850
rect 96682 65798 100832 65850
rect 1104 65776 100832 65798
rect 1104 65306 100832 65328
rect 1104 65254 4874 65306
rect 4926 65254 4938 65306
rect 4990 65254 5002 65306
rect 5054 65254 5066 65306
rect 5118 65254 5130 65306
rect 5182 65254 35594 65306
rect 35646 65254 35658 65306
rect 35710 65254 35722 65306
rect 35774 65254 35786 65306
rect 35838 65254 35850 65306
rect 35902 65254 66314 65306
rect 66366 65254 66378 65306
rect 66430 65254 66442 65306
rect 66494 65254 66506 65306
rect 66558 65254 66570 65306
rect 66622 65254 97034 65306
rect 97086 65254 97098 65306
rect 97150 65254 97162 65306
rect 97214 65254 97226 65306
rect 97278 65254 97290 65306
rect 97342 65254 100832 65306
rect 1104 65232 100832 65254
rect 1104 64762 100832 64784
rect 1104 64710 4214 64762
rect 4266 64710 4278 64762
rect 4330 64710 4342 64762
rect 4394 64710 4406 64762
rect 4458 64710 4470 64762
rect 4522 64710 34934 64762
rect 34986 64710 34998 64762
rect 35050 64710 35062 64762
rect 35114 64710 35126 64762
rect 35178 64710 35190 64762
rect 35242 64710 65654 64762
rect 65706 64710 65718 64762
rect 65770 64710 65782 64762
rect 65834 64710 65846 64762
rect 65898 64710 65910 64762
rect 65962 64710 96374 64762
rect 96426 64710 96438 64762
rect 96490 64710 96502 64762
rect 96554 64710 96566 64762
rect 96618 64710 96630 64762
rect 96682 64710 100832 64762
rect 1104 64688 100832 64710
rect 1104 64218 100832 64240
rect 1104 64166 4874 64218
rect 4926 64166 4938 64218
rect 4990 64166 5002 64218
rect 5054 64166 5066 64218
rect 5118 64166 5130 64218
rect 5182 64166 35594 64218
rect 35646 64166 35658 64218
rect 35710 64166 35722 64218
rect 35774 64166 35786 64218
rect 35838 64166 35850 64218
rect 35902 64166 66314 64218
rect 66366 64166 66378 64218
rect 66430 64166 66442 64218
rect 66494 64166 66506 64218
rect 66558 64166 66570 64218
rect 66622 64166 97034 64218
rect 97086 64166 97098 64218
rect 97150 64166 97162 64218
rect 97214 64166 97226 64218
rect 97278 64166 97290 64218
rect 97342 64166 100832 64218
rect 1104 64144 100832 64166
rect 1104 63674 100832 63696
rect 1104 63622 4214 63674
rect 4266 63622 4278 63674
rect 4330 63622 4342 63674
rect 4394 63622 4406 63674
rect 4458 63622 4470 63674
rect 4522 63622 34934 63674
rect 34986 63622 34998 63674
rect 35050 63622 35062 63674
rect 35114 63622 35126 63674
rect 35178 63622 35190 63674
rect 35242 63622 65654 63674
rect 65706 63622 65718 63674
rect 65770 63622 65782 63674
rect 65834 63622 65846 63674
rect 65898 63622 65910 63674
rect 65962 63622 96374 63674
rect 96426 63622 96438 63674
rect 96490 63622 96502 63674
rect 96554 63622 96566 63674
rect 96618 63622 96630 63674
rect 96682 63622 100832 63674
rect 1104 63600 100832 63622
rect 1104 63130 100832 63152
rect 1104 63078 4874 63130
rect 4926 63078 4938 63130
rect 4990 63078 5002 63130
rect 5054 63078 5066 63130
rect 5118 63078 5130 63130
rect 5182 63078 35594 63130
rect 35646 63078 35658 63130
rect 35710 63078 35722 63130
rect 35774 63078 35786 63130
rect 35838 63078 35850 63130
rect 35902 63078 66314 63130
rect 66366 63078 66378 63130
rect 66430 63078 66442 63130
rect 66494 63078 66506 63130
rect 66558 63078 66570 63130
rect 66622 63078 97034 63130
rect 97086 63078 97098 63130
rect 97150 63078 97162 63130
rect 97214 63078 97226 63130
rect 97278 63078 97290 63130
rect 97342 63078 100832 63130
rect 1104 63056 100832 63078
rect 96246 62840 96252 62892
rect 96304 62880 96310 62892
rect 100205 62883 100263 62889
rect 100205 62880 100217 62883
rect 96304 62852 100217 62880
rect 96304 62840 96310 62852
rect 100205 62849 100217 62852
rect 100251 62849 100263 62883
rect 100205 62843 100263 62849
rect 100386 62636 100392 62688
rect 100444 62636 100450 62688
rect 1104 62586 100832 62608
rect 1104 62534 4214 62586
rect 4266 62534 4278 62586
rect 4330 62534 4342 62586
rect 4394 62534 4406 62586
rect 4458 62534 4470 62586
rect 4522 62534 34934 62586
rect 34986 62534 34998 62586
rect 35050 62534 35062 62586
rect 35114 62534 35126 62586
rect 35178 62534 35190 62586
rect 35242 62534 65654 62586
rect 65706 62534 65718 62586
rect 65770 62534 65782 62586
rect 65834 62534 65846 62586
rect 65898 62534 65910 62586
rect 65962 62534 96374 62586
rect 96426 62534 96438 62586
rect 96490 62534 96502 62586
rect 96554 62534 96566 62586
rect 96618 62534 96630 62586
rect 96682 62534 100832 62586
rect 1104 62512 100832 62534
rect 1673 62271 1731 62277
rect 1673 62237 1685 62271
rect 1719 62268 1731 62271
rect 1719 62240 1900 62268
rect 1719 62237 1731 62240
rect 1673 62231 1731 62237
rect 1872 62144 1900 62240
rect 96890 62228 96896 62280
rect 96948 62268 96954 62280
rect 100205 62271 100263 62277
rect 100205 62268 100217 62271
rect 96948 62240 100217 62268
rect 96948 62228 96954 62240
rect 100205 62237 100217 62240
rect 100251 62237 100263 62271
rect 100205 62231 100263 62237
rect 1486 62092 1492 62144
rect 1544 62092 1550 62144
rect 1854 62092 1860 62144
rect 1912 62092 1918 62144
rect 100386 62092 100392 62144
rect 100444 62092 100450 62144
rect 1104 62042 100832 62064
rect 1104 61990 4874 62042
rect 4926 61990 4938 62042
rect 4990 61990 5002 62042
rect 5054 61990 5066 62042
rect 5118 61990 5130 62042
rect 5182 61990 35594 62042
rect 35646 61990 35658 62042
rect 35710 61990 35722 62042
rect 35774 61990 35786 62042
rect 35838 61990 35850 62042
rect 35902 61990 66314 62042
rect 66366 61990 66378 62042
rect 66430 61990 66442 62042
rect 66494 61990 66506 62042
rect 66558 61990 66570 62042
rect 66622 61990 97034 62042
rect 97086 61990 97098 62042
rect 97150 61990 97162 62042
rect 97214 61990 97226 62042
rect 97278 61990 97290 62042
rect 97342 61990 100832 62042
rect 1104 61968 100832 61990
rect 1673 61795 1731 61801
rect 1673 61761 1685 61795
rect 1719 61792 1731 61795
rect 21082 61792 21088 61804
rect 1719 61764 21088 61792
rect 1719 61761 1731 61764
rect 1673 61755 1731 61761
rect 21082 61752 21088 61764
rect 21140 61752 21146 61804
rect 100202 61752 100208 61804
rect 100260 61752 100266 61804
rect 842 61548 848 61600
rect 900 61588 906 61600
rect 1489 61591 1547 61597
rect 1489 61588 1501 61591
rect 900 61560 1501 61588
rect 900 61548 906 61560
rect 1489 61557 1501 61560
rect 1535 61557 1547 61591
rect 1489 61551 1547 61557
rect 100386 61548 100392 61600
rect 100444 61548 100450 61600
rect 1104 61498 100832 61520
rect 1104 61446 4214 61498
rect 4266 61446 4278 61498
rect 4330 61446 4342 61498
rect 4394 61446 4406 61498
rect 4458 61446 4470 61498
rect 4522 61446 34934 61498
rect 34986 61446 34998 61498
rect 35050 61446 35062 61498
rect 35114 61446 35126 61498
rect 35178 61446 35190 61498
rect 35242 61446 65654 61498
rect 65706 61446 65718 61498
rect 65770 61446 65782 61498
rect 65834 61446 65846 61498
rect 65898 61446 65910 61498
rect 65962 61446 96374 61498
rect 96426 61446 96438 61498
rect 96490 61446 96502 61498
rect 96554 61446 96566 61498
rect 96618 61446 96630 61498
rect 96682 61446 100832 61498
rect 1104 61424 100832 61446
rect 21082 61344 21088 61396
rect 21140 61344 21146 61396
rect 77110 61344 77116 61396
rect 77168 61384 77174 61396
rect 81897 61387 81955 61393
rect 81897 61384 81909 61387
rect 77168 61356 81909 61384
rect 77168 61344 77174 61356
rect 81897 61353 81909 61356
rect 81943 61384 81955 61387
rect 82338 61387 82396 61393
rect 82338 61384 82350 61387
rect 81943 61356 82350 61384
rect 81943 61353 81955 61356
rect 81897 61347 81955 61353
rect 82338 61353 82350 61356
rect 82384 61353 82396 61387
rect 82338 61347 82396 61353
rect 82446 61344 82452 61396
rect 82504 61384 82510 61396
rect 96246 61384 96252 61396
rect 82504 61356 96252 61384
rect 82504 61344 82510 61356
rect 96246 61344 96252 61356
rect 96304 61344 96310 61396
rect 22557 61251 22615 61257
rect 22557 61217 22569 61251
rect 22603 61248 22615 61251
rect 28166 61248 28172 61260
rect 22603 61220 28172 61248
rect 22603 61217 22615 61220
rect 22557 61211 22615 61217
rect 28166 61208 28172 61220
rect 28224 61208 28230 61260
rect 78861 61251 78919 61257
rect 78861 61248 78873 61251
rect 77036 61220 78873 61248
rect 77036 61192 77064 61220
rect 78861 61217 78873 61220
rect 78907 61248 78919 61251
rect 79686 61248 79692 61260
rect 78907 61220 79692 61248
rect 78907 61217 78919 61220
rect 78861 61211 78919 61217
rect 79686 61208 79692 61220
rect 79744 61208 79750 61260
rect 79870 61208 79876 61260
rect 79928 61248 79934 61260
rect 80609 61251 80667 61257
rect 79928 61220 80376 61248
rect 79928 61208 79934 61220
rect 22830 61140 22836 61192
rect 22888 61140 22894 61192
rect 77018 61140 77024 61192
rect 77076 61140 77082 61192
rect 80348 61180 80376 61220
rect 80609 61217 80621 61251
rect 80655 61248 80667 61251
rect 96890 61248 96896 61260
rect 80655 61220 96896 61248
rect 80655 61217 80667 61220
rect 80609 61211 80667 61217
rect 96890 61208 96896 61220
rect 96948 61208 96954 61260
rect 80701 61183 80759 61189
rect 80701 61180 80713 61183
rect 80348 61152 80713 61180
rect 80701 61149 80713 61152
rect 80747 61149 80759 61183
rect 80701 61143 80759 61149
rect 81526 61140 81532 61192
rect 81584 61180 81590 61192
rect 82081 61183 82139 61189
rect 82081 61180 82093 61183
rect 81584 61152 82093 61180
rect 81584 61140 81590 61152
rect 82081 61149 82093 61152
rect 82127 61149 82139 61183
rect 82081 61143 82139 61149
rect 83918 61140 83924 61192
rect 83976 61140 83982 61192
rect 77297 61115 77355 61121
rect 22126 61084 24440 61112
rect 24412 61044 24440 61084
rect 77297 61081 77309 61115
rect 77343 61081 77355 61115
rect 77297 61075 77355 61081
rect 28810 61044 28816 61056
rect 24412 61016 28816 61044
rect 28810 61004 28816 61016
rect 28868 61004 28874 61056
rect 71774 61004 71780 61056
rect 71832 61044 71838 61056
rect 76837 61047 76895 61053
rect 76837 61044 76849 61047
rect 71832 61016 76849 61044
rect 71832 61004 71838 61016
rect 76837 61013 76849 61016
rect 76883 61044 76895 61047
rect 77312 61044 77340 61075
rect 77754 61072 77760 61124
rect 77812 61072 77818 61124
rect 79134 61072 79140 61124
rect 79192 61072 79198 61124
rect 79594 61072 79600 61124
rect 79652 61072 79658 61124
rect 82446 61112 82452 61124
rect 80624 61084 82452 61112
rect 76883 61016 77340 61044
rect 78769 61047 78827 61053
rect 76883 61013 76895 61016
rect 76837 61007 76895 61013
rect 78769 61013 78781 61047
rect 78815 61044 78827 61047
rect 80624 61044 80652 61084
rect 82446 61072 82452 61084
rect 82504 61072 82510 61124
rect 82814 61072 82820 61124
rect 82872 61072 82878 61124
rect 78815 61016 80652 61044
rect 78815 61013 78827 61016
rect 78769 61007 78827 61013
rect 83826 61004 83832 61056
rect 83884 61004 83890 61056
rect 84010 61004 84016 61056
rect 84068 61004 84074 61056
rect 1104 60954 100832 60976
rect 1104 60902 4874 60954
rect 4926 60902 4938 60954
rect 4990 60902 5002 60954
rect 5054 60902 5066 60954
rect 5118 60902 5130 60954
rect 5182 60902 35594 60954
rect 35646 60902 35658 60954
rect 35710 60902 35722 60954
rect 35774 60902 35786 60954
rect 35838 60902 35850 60954
rect 35902 60902 66314 60954
rect 66366 60902 66378 60954
rect 66430 60902 66442 60954
rect 66494 60902 66506 60954
rect 66558 60902 66570 60954
rect 66622 60902 97034 60954
rect 97086 60902 97098 60954
rect 97150 60902 97162 60954
rect 97214 60902 97226 60954
rect 97278 60902 97290 60954
rect 97342 60902 100832 60954
rect 1104 60880 100832 60902
rect 30377 60843 30435 60849
rect 30377 60840 30389 60843
rect 24228 60812 30389 60840
rect 24228 60772 24256 60812
rect 30377 60809 30389 60812
rect 30423 60809 30435 60843
rect 30377 60803 30435 60809
rect 79134 60800 79140 60852
rect 79192 60840 79198 60852
rect 79870 60840 79876 60852
rect 79192 60812 79876 60840
rect 79192 60800 79198 60812
rect 79870 60800 79876 60812
rect 79928 60800 79934 60852
rect 83826 60800 83832 60852
rect 83884 60840 83890 60852
rect 83884 60812 100248 60840
rect 83884 60800 83890 60812
rect 48133 60775 48191 60781
rect 48133 60772 48145 60775
rect 23598 60744 24256 60772
rect 24320 60744 48145 60772
rect 24026 60596 24032 60648
rect 24084 60596 24090 60648
rect 24320 60645 24348 60744
rect 48133 60741 48145 60744
rect 48179 60772 48191 60775
rect 48406 60772 48412 60784
rect 48179 60744 48412 60772
rect 48179 60741 48191 60744
rect 48133 60735 48191 60741
rect 48406 60732 48412 60744
rect 48464 60772 48470 60784
rect 49418 60772 49424 60784
rect 48464 60744 49424 60772
rect 48464 60732 48470 60744
rect 49418 60732 49424 60744
rect 49476 60732 49482 60784
rect 79612 60744 80454 60772
rect 28810 60664 28816 60716
rect 28868 60704 28874 60716
rect 29181 60707 29239 60713
rect 29181 60704 29193 60707
rect 28868 60676 29193 60704
rect 28868 60664 28874 60676
rect 29181 60673 29193 60676
rect 29227 60673 29239 60707
rect 29181 60667 29239 60673
rect 29273 60707 29331 60713
rect 29273 60673 29285 60707
rect 29319 60704 29331 60707
rect 30469 60707 30527 60713
rect 30469 60704 30481 60707
rect 29319 60676 30481 60704
rect 29319 60673 29331 60676
rect 29273 60667 29331 60673
rect 30469 60673 30481 60676
rect 30515 60704 30527 60707
rect 46658 60704 46664 60716
rect 30515 60676 46664 60704
rect 30515 60673 30527 60676
rect 30469 60667 30527 60673
rect 46658 60664 46664 60676
rect 46716 60664 46722 60716
rect 77205 60707 77263 60713
rect 77205 60673 77217 60707
rect 77251 60704 77263 60707
rect 78493 60707 78551 60713
rect 78493 60704 78505 60707
rect 77251 60676 78505 60704
rect 77251 60673 77263 60676
rect 77205 60667 77263 60673
rect 78493 60673 78505 60676
rect 78539 60704 78551 60707
rect 79226 60704 79232 60716
rect 78539 60676 79232 60704
rect 78539 60673 78551 60676
rect 78493 60667 78551 60673
rect 79226 60664 79232 60676
rect 79284 60664 79290 60716
rect 79321 60707 79379 60713
rect 79321 60673 79333 60707
rect 79367 60704 79379 60707
rect 79612 60704 79640 60744
rect 81710 60732 81716 60784
rect 81768 60772 81774 60784
rect 81768 60744 82294 60772
rect 81768 60732 81774 60744
rect 84010 60732 84016 60784
rect 84068 60772 84074 60784
rect 84068 60744 84502 60772
rect 84068 60732 84074 60744
rect 85574 60732 85580 60784
rect 85632 60772 85638 60784
rect 85632 60744 86434 60772
rect 85632 60732 85638 60744
rect 79367 60676 79640 60704
rect 79367 60673 79379 60676
rect 79321 60667 79379 60673
rect 79686 60664 79692 60716
rect 79744 60664 79750 60716
rect 100220 60713 100248 60812
rect 100205 60707 100263 60713
rect 100205 60673 100217 60707
rect 100251 60673 100263 60707
rect 100205 60667 100263 60673
rect 24305 60639 24363 60645
rect 24305 60636 24317 60639
rect 24228 60608 24317 60636
rect 22557 60571 22615 60577
rect 22557 60568 22569 60571
rect 6886 60540 22569 60568
rect 1854 60460 1860 60512
rect 1912 60500 1918 60512
rect 6886 60500 6914 60540
rect 22557 60537 22569 60540
rect 22603 60537 22615 60571
rect 22557 60531 22615 60537
rect 1912 60472 6914 60500
rect 1912 60460 1918 60472
rect 22370 60460 22376 60512
rect 22428 60500 22434 60512
rect 22830 60500 22836 60512
rect 22428 60472 22836 60500
rect 22428 60460 22434 60472
rect 22830 60460 22836 60472
rect 22888 60500 22894 60512
rect 24228 60500 24256 60608
rect 24305 60605 24317 60608
rect 24351 60605 24363 60639
rect 24305 60599 24363 60605
rect 77113 60639 77171 60645
rect 77113 60605 77125 60639
rect 77159 60636 77171 60639
rect 77754 60636 77760 60648
rect 77159 60608 77760 60636
rect 77159 60605 77171 60608
rect 77113 60599 77171 60605
rect 77754 60596 77760 60608
rect 77812 60596 77818 60648
rect 78585 60639 78643 60645
rect 78585 60605 78597 60639
rect 78631 60636 78643 60639
rect 79594 60636 79600 60648
rect 78631 60608 79600 60636
rect 78631 60605 78643 60608
rect 78585 60599 78643 60605
rect 79594 60596 79600 60608
rect 79652 60596 79658 60648
rect 79965 60639 80023 60645
rect 79965 60636 79977 60639
rect 79704 60608 79977 60636
rect 79704 60568 79732 60608
rect 79965 60605 79977 60608
rect 80011 60605 80023 60639
rect 79965 60599 80023 60605
rect 81526 60596 81532 60648
rect 81584 60596 81590 60648
rect 81802 60596 81808 60648
rect 81860 60636 81866 60648
rect 83369 60639 83427 60645
rect 83369 60636 83381 60639
rect 81860 60608 83381 60636
rect 81860 60596 81866 60608
rect 83369 60605 83381 60608
rect 83415 60605 83427 60639
rect 83369 60599 83427 60605
rect 83918 60596 83924 60648
rect 83976 60596 83982 60648
rect 85666 60596 85672 60648
rect 85724 60596 85730 60648
rect 85945 60639 86003 60645
rect 85945 60605 85957 60639
rect 85991 60636 86003 60639
rect 85991 60608 86264 60636
rect 85991 60605 86003 60608
rect 85945 60599 86003 60605
rect 81544 60568 81572 60596
rect 79520 60540 79732 60568
rect 81360 60540 81572 60568
rect 79520 60512 79548 60540
rect 22888 60472 24256 60500
rect 22888 60460 22894 60472
rect 79502 60460 79508 60512
rect 79560 60460 79566 60512
rect 79686 60460 79692 60512
rect 79744 60500 79750 60512
rect 81360 60500 81388 60540
rect 79744 60472 81388 60500
rect 79744 60460 79750 60472
rect 81434 60460 81440 60512
rect 81492 60460 81498 60512
rect 81544 60500 81572 60540
rect 82832 60540 83504 60568
rect 82832 60500 82860 60540
rect 81544 60472 82860 60500
rect 83274 60460 83280 60512
rect 83332 60460 83338 60512
rect 83476 60500 83504 60540
rect 85960 60500 85988 60599
rect 83476 60472 85988 60500
rect 86126 60460 86132 60512
rect 86184 60460 86190 60512
rect 86236 60500 86264 60608
rect 87598 60596 87604 60648
rect 87656 60596 87662 60648
rect 87874 60596 87880 60648
rect 87932 60596 87938 60648
rect 100386 60528 100392 60580
rect 100444 60528 100450 60580
rect 87874 60500 87880 60512
rect 86236 60472 87880 60500
rect 87874 60460 87880 60472
rect 87932 60460 87938 60512
rect 1104 60410 100832 60432
rect 1104 60358 1322 60410
rect 1374 60358 1386 60410
rect 1438 60358 4214 60410
rect 4266 60358 4278 60410
rect 4330 60358 4342 60410
rect 4394 60358 4406 60410
rect 4458 60358 4470 60410
rect 4522 60358 34934 60410
rect 34986 60358 34998 60410
rect 35050 60358 35062 60410
rect 35114 60358 35126 60410
rect 35178 60358 35190 60410
rect 35242 60358 65654 60410
rect 65706 60358 65718 60410
rect 65770 60358 65782 60410
rect 65834 60358 65846 60410
rect 65898 60358 65910 60410
rect 65962 60358 96374 60410
rect 96426 60358 96438 60410
rect 96490 60358 96502 60410
rect 96554 60358 96566 60410
rect 96618 60358 96630 60410
rect 96682 60358 98930 60410
rect 98982 60358 98994 60410
rect 99046 60358 99058 60410
rect 99110 60358 99122 60410
rect 99174 60358 99186 60410
rect 99238 60358 100832 60410
rect 1104 60336 100832 60358
rect 24026 60256 24032 60308
rect 24084 60296 24090 60308
rect 29178 60296 29184 60308
rect 24084 60268 29184 60296
rect 24084 60256 24090 60268
rect 29178 60256 29184 60268
rect 29236 60256 29242 60308
rect 48406 60256 48412 60308
rect 48464 60256 48470 60308
rect 80241 60299 80299 60305
rect 80241 60265 80253 60299
rect 80287 60296 80299 60299
rect 81710 60296 81716 60308
rect 80287 60268 81716 60296
rect 80287 60265 80299 60268
rect 80241 60259 80299 60265
rect 81710 60256 81716 60268
rect 81768 60256 81774 60308
rect 81805 60299 81863 60305
rect 81805 60265 81817 60299
rect 81851 60296 81863 60299
rect 82814 60296 82820 60308
rect 81851 60268 82820 60296
rect 81851 60265 81863 60268
rect 81805 60259 81863 60265
rect 82814 60256 82820 60268
rect 82872 60256 82878 60308
rect 84473 60299 84531 60305
rect 84473 60265 84485 60299
rect 84519 60296 84531 60299
rect 85574 60296 85580 60308
rect 84519 60268 85580 60296
rect 84519 60265 84531 60268
rect 84473 60259 84531 60265
rect 85574 60256 85580 60268
rect 85632 60256 85638 60308
rect 85666 60256 85672 60308
rect 85724 60296 85730 60308
rect 85945 60299 86003 60305
rect 85945 60296 85957 60299
rect 85724 60268 85957 60296
rect 85724 60256 85730 60268
rect 85945 60265 85957 60268
rect 85991 60265 86003 60299
rect 85945 60259 86003 60265
rect 87598 60256 87604 60308
rect 87656 60296 87662 60308
rect 87693 60299 87751 60305
rect 87693 60296 87705 60299
rect 87656 60268 87705 60296
rect 87656 60256 87662 60268
rect 87693 60265 87705 60268
rect 87739 60265 87751 60299
rect 100202 60296 100208 60308
rect 87693 60259 87751 60265
rect 89686 60268 100208 60296
rect 83274 60188 83280 60240
rect 83332 60228 83338 60240
rect 89686 60228 89714 60268
rect 100202 60256 100208 60268
rect 100260 60256 100266 60308
rect 83332 60200 89714 60228
rect 83332 60188 83338 60200
rect 91738 60188 91744 60240
rect 91796 60228 91802 60240
rect 91796 60200 100248 60228
rect 91796 60188 91802 60200
rect 75457 60163 75515 60169
rect 75457 60129 75469 60163
rect 75503 60160 75515 60163
rect 77018 60160 77024 60172
rect 75503 60132 77024 60160
rect 75503 60129 75515 60132
rect 75457 60123 75515 60129
rect 77018 60120 77024 60132
rect 77076 60120 77082 60172
rect 83918 60120 83924 60172
rect 83976 60160 83982 60172
rect 85117 60163 85175 60169
rect 85117 60160 85129 60163
rect 83976 60132 85129 60160
rect 83976 60120 83982 60132
rect 85117 60129 85129 60132
rect 85163 60160 85175 60163
rect 87601 60163 87659 60169
rect 85163 60132 87552 60160
rect 85163 60129 85175 60132
rect 85117 60123 85175 60129
rect 79226 60052 79232 60104
rect 79284 60092 79290 60104
rect 80149 60095 80207 60101
rect 80149 60092 80161 60095
rect 79284 60064 80161 60092
rect 79284 60052 79290 60064
rect 80149 60061 80161 60064
rect 80195 60092 80207 60095
rect 81342 60092 81348 60104
rect 80195 60064 81348 60092
rect 80195 60061 80207 60064
rect 80149 60055 80207 60061
rect 81342 60052 81348 60064
rect 81400 60052 81406 60104
rect 81713 60095 81771 60101
rect 81713 60061 81725 60095
rect 81759 60092 81771 60095
rect 83826 60092 83832 60104
rect 81759 60064 83832 60092
rect 81759 60061 81771 60064
rect 81713 60055 81771 60061
rect 83826 60052 83832 60064
rect 83884 60092 83890 60104
rect 84378 60092 84384 60104
rect 83884 60064 84384 60092
rect 83884 60052 83890 60064
rect 84378 60052 84384 60064
rect 84436 60052 84442 60104
rect 85761 60095 85819 60101
rect 85761 60061 85773 60095
rect 85807 60092 85819 60095
rect 85853 60095 85911 60101
rect 85853 60092 85865 60095
rect 85807 60064 85865 60092
rect 85807 60061 85819 60064
rect 85761 60055 85819 60061
rect 85853 60061 85865 60064
rect 85899 60061 85911 60095
rect 85853 60055 85911 60061
rect 86126 60052 86132 60104
rect 86184 60092 86190 60104
rect 86957 60095 87015 60101
rect 86957 60092 86969 60095
rect 86184 60064 86969 60092
rect 86184 60052 86190 60064
rect 86957 60061 86969 60064
rect 87003 60061 87015 60095
rect 87524 60092 87552 60132
rect 87601 60129 87613 60163
rect 87647 60160 87659 60163
rect 87969 60163 88027 60169
rect 87969 60160 87981 60163
rect 87647 60132 87981 60160
rect 87647 60129 87659 60132
rect 87601 60123 87659 60129
rect 87969 60129 87981 60132
rect 88015 60129 88027 60163
rect 87969 60123 88027 60129
rect 88061 60095 88119 60101
rect 88061 60092 88073 60095
rect 87524 60064 88073 60092
rect 86957 60055 87015 60061
rect 88061 60061 88073 60064
rect 88107 60092 88119 60095
rect 89530 60092 89536 60104
rect 88107 60064 89536 60092
rect 88107 60061 88119 60064
rect 88061 60055 88119 60061
rect 89530 60052 89536 60064
rect 89588 60052 89594 60104
rect 89714 60052 89720 60104
rect 89772 60092 89778 60104
rect 98362 60092 98368 60104
rect 89772 60064 98368 60092
rect 89772 60052 89778 60064
rect 98362 60052 98368 60064
rect 98420 60052 98426 60104
rect 100220 60101 100248 60200
rect 100205 60095 100263 60101
rect 100205 60061 100217 60095
rect 100251 60061 100263 60095
rect 100205 60055 100263 60061
rect 49881 60027 49939 60033
rect 49881 59993 49893 60027
rect 49927 60024 49939 60027
rect 49927 59996 55214 60024
rect 49927 59993 49939 59996
rect 49881 59987 49939 59993
rect 55186 59956 55214 59996
rect 57054 59984 57060 60036
rect 57112 59984 57118 60036
rect 73709 60027 73767 60033
rect 73709 60024 73721 60027
rect 64846 59996 73721 60024
rect 55769 59959 55827 59965
rect 55769 59956 55781 59959
rect 55186 59928 55781 59956
rect 55769 59925 55781 59928
rect 55815 59956 55827 59959
rect 64846 59956 64874 59996
rect 73709 59993 73721 59996
rect 73755 59993 73767 60027
rect 73709 59987 73767 59993
rect 81434 59984 81440 60036
rect 81492 60024 81498 60036
rect 91738 60024 91744 60036
rect 81492 59996 91744 60024
rect 81492 59984 81498 59996
rect 91738 59984 91744 59996
rect 91796 59984 91802 60036
rect 55815 59928 64874 59956
rect 55815 59925 55827 59928
rect 55769 59919 55827 59925
rect 100386 59916 100392 59968
rect 100444 59916 100450 59968
rect 1104 59866 100832 59888
rect 1104 59814 1690 59866
rect 1742 59814 1754 59866
rect 1806 59814 4874 59866
rect 4926 59814 4938 59866
rect 4990 59814 5002 59866
rect 5054 59814 5066 59866
rect 5118 59814 5130 59866
rect 5182 59814 35594 59866
rect 35646 59814 35658 59866
rect 35710 59814 35722 59866
rect 35774 59814 35786 59866
rect 35838 59814 35850 59866
rect 35902 59814 66314 59866
rect 66366 59814 66378 59866
rect 66430 59814 66442 59866
rect 66494 59814 66506 59866
rect 66558 59814 66570 59866
rect 66622 59814 97034 59866
rect 97086 59814 97098 59866
rect 97150 59814 97162 59866
rect 97214 59814 97226 59866
rect 97278 59814 97290 59866
rect 97342 59814 99666 59866
rect 99718 59814 99730 59866
rect 99782 59814 99794 59866
rect 99846 59814 99858 59866
rect 99910 59814 99922 59866
rect 99974 59814 100832 59866
rect 1104 59792 100832 59814
rect 2682 59372 2688 59424
rect 2740 59412 2746 59424
rect 22370 59412 22376 59424
rect 2740 59384 22376 59412
rect 2740 59372 2746 59384
rect 22370 59372 22376 59384
rect 22428 59372 22434 59424
rect 1104 59322 1932 59344
rect 1104 59270 1322 59322
rect 1374 59270 1386 59322
rect 1438 59270 1932 59322
rect 1104 59248 1932 59270
rect 97980 59322 100832 59344
rect 97980 59270 98930 59322
rect 98982 59270 98994 59322
rect 99046 59270 99058 59322
rect 99110 59270 99122 59322
rect 99174 59270 99186 59322
rect 99238 59270 100832 59322
rect 97980 59248 100832 59270
rect 1104 58778 1932 58800
rect 1104 58726 1690 58778
rect 1742 58726 1754 58778
rect 1806 58726 1932 58778
rect 84378 58760 84384 58812
rect 84436 58800 84442 58812
rect 97350 58800 97356 58812
rect 84436 58772 97356 58800
rect 84436 58760 84442 58772
rect 97350 58760 97356 58772
rect 97408 58760 97414 58812
rect 97980 58778 100832 58800
rect 1104 58704 1932 58726
rect 81342 58692 81348 58744
rect 81400 58732 81406 58744
rect 97442 58732 97448 58744
rect 81400 58704 97448 58732
rect 81400 58692 81406 58704
rect 97442 58692 97448 58704
rect 97500 58692 97506 58744
rect 97980 58726 99666 58778
rect 99718 58726 99730 58778
rect 99782 58726 99794 58778
rect 99846 58726 99858 58778
rect 99910 58726 99922 58778
rect 99974 58726 100832 58778
rect 97980 58704 100832 58726
rect 57054 58624 57060 58676
rect 57112 58664 57118 58676
rect 97258 58664 97264 58676
rect 57112 58636 97264 58664
rect 57112 58624 57118 58636
rect 97258 58624 97264 58636
rect 97316 58624 97322 58676
rect 1104 58234 1932 58256
rect 1104 58182 1322 58234
rect 1374 58182 1386 58234
rect 1438 58182 1932 58234
rect 1104 58160 1932 58182
rect 97980 58234 100832 58256
rect 97980 58182 98930 58234
rect 98982 58182 98994 58234
rect 99046 58182 99058 58234
rect 99110 58182 99122 58234
rect 99174 58182 99186 58234
rect 99238 58182 100832 58234
rect 97980 58160 100832 58182
rect 1104 57690 1932 57712
rect 1104 57638 1690 57690
rect 1742 57638 1754 57690
rect 1806 57638 1932 57690
rect 1104 57616 1932 57638
rect 97980 57690 100832 57712
rect 97980 57638 99666 57690
rect 99718 57638 99730 57690
rect 99782 57638 99794 57690
rect 99846 57638 99858 57690
rect 99910 57638 99922 57690
rect 99974 57638 100832 57690
rect 97980 57616 100832 57638
rect 1104 57146 1932 57168
rect 1104 57094 1322 57146
rect 1374 57094 1386 57146
rect 1438 57094 1932 57146
rect 1104 57072 1932 57094
rect 97980 57146 100832 57168
rect 97980 57094 98930 57146
rect 98982 57094 98994 57146
rect 99046 57094 99058 57146
rect 99110 57094 99122 57146
rect 99174 57094 99186 57146
rect 99238 57094 100832 57146
rect 97980 57072 100832 57094
rect 1104 56602 1932 56624
rect 1104 56550 1690 56602
rect 1742 56550 1754 56602
rect 1806 56550 1932 56602
rect 1104 56528 1932 56550
rect 97980 56602 100832 56624
rect 97980 56550 99666 56602
rect 99718 56550 99730 56602
rect 99782 56550 99794 56602
rect 99846 56550 99858 56602
rect 99910 56550 99922 56602
rect 99974 56550 100832 56602
rect 97980 56528 100832 56550
rect 1104 56058 1932 56080
rect 1104 56006 1322 56058
rect 1374 56006 1386 56058
rect 1438 56006 1932 56058
rect 1104 55984 1932 56006
rect 97980 56058 100832 56080
rect 97980 56006 98930 56058
rect 98982 56006 98994 56058
rect 99046 56006 99058 56058
rect 99110 56006 99122 56058
rect 99174 56006 99186 56058
rect 99238 56006 100832 56058
rect 97980 55984 100832 56006
rect 1104 55514 1932 55536
rect 1104 55462 1690 55514
rect 1742 55462 1754 55514
rect 1806 55462 1932 55514
rect 1104 55440 1932 55462
rect 97980 55514 100832 55536
rect 97980 55462 99666 55514
rect 99718 55462 99730 55514
rect 99782 55462 99794 55514
rect 99846 55462 99858 55514
rect 99910 55462 99922 55514
rect 99974 55462 100832 55514
rect 97980 55440 100832 55462
rect 1104 54970 1932 54992
rect 1104 54918 1322 54970
rect 1374 54918 1386 54970
rect 1438 54918 1932 54970
rect 1104 54896 1932 54918
rect 97980 54970 100832 54992
rect 97980 54918 98930 54970
rect 98982 54918 98994 54970
rect 99046 54918 99058 54970
rect 99110 54918 99122 54970
rect 99174 54918 99186 54970
rect 99238 54918 100832 54970
rect 97980 54896 100832 54918
rect 1104 54426 1932 54448
rect 1104 54374 1690 54426
rect 1742 54374 1754 54426
rect 1806 54374 1932 54426
rect 1104 54352 1932 54374
rect 97980 54426 100832 54448
rect 97980 54374 99666 54426
rect 99718 54374 99730 54426
rect 99782 54374 99794 54426
rect 99846 54374 99858 54426
rect 99910 54374 99922 54426
rect 99974 54374 100832 54426
rect 97980 54352 100832 54374
rect 97074 53932 97080 53984
rect 97132 53972 97138 53984
rect 98273 53975 98331 53981
rect 98273 53972 98285 53975
rect 97132 53944 98285 53972
rect 97132 53932 97138 53944
rect 98273 53941 98285 53944
rect 98319 53941 98331 53975
rect 98273 53935 98331 53941
rect 1104 53882 1932 53904
rect 1104 53830 1322 53882
rect 1374 53830 1386 53882
rect 1438 53830 1932 53882
rect 1104 53808 1932 53830
rect 97980 53882 100832 53904
rect 97980 53830 98930 53882
rect 98982 53830 98994 53882
rect 99046 53830 99058 53882
rect 99110 53830 99122 53882
rect 99174 53830 99186 53882
rect 99238 53830 100832 53882
rect 97980 53808 100832 53830
rect 1104 53338 1932 53360
rect 1104 53286 1690 53338
rect 1742 53286 1754 53338
rect 1806 53286 1932 53338
rect 1104 53264 1932 53286
rect 97980 53338 100832 53360
rect 97980 53286 99666 53338
rect 99718 53286 99730 53338
rect 99782 53286 99794 53338
rect 99846 53286 99858 53338
rect 99910 53286 99922 53338
rect 99974 53286 100832 53338
rect 97980 53264 100832 53286
rect 1104 52794 1932 52816
rect 1104 52742 1322 52794
rect 1374 52742 1386 52794
rect 1438 52742 1932 52794
rect 1104 52720 1932 52742
rect 97980 52794 100832 52816
rect 97980 52742 98930 52794
rect 98982 52742 98994 52794
rect 99046 52742 99058 52794
rect 99110 52742 99122 52794
rect 99174 52742 99186 52794
rect 99238 52742 100832 52794
rect 97980 52720 100832 52742
rect 1104 52250 1932 52272
rect 1104 52198 1690 52250
rect 1742 52198 1754 52250
rect 1806 52198 1932 52250
rect 1104 52176 1932 52198
rect 97980 52250 100832 52272
rect 97980 52198 99666 52250
rect 99718 52198 99730 52250
rect 99782 52198 99794 52250
rect 99846 52198 99858 52250
rect 99910 52198 99922 52250
rect 99974 52198 100832 52250
rect 97980 52176 100832 52198
rect 1104 51706 1932 51728
rect 1104 51654 1322 51706
rect 1374 51654 1386 51706
rect 1438 51654 1932 51706
rect 1104 51632 1932 51654
rect 97980 51706 100832 51728
rect 97980 51654 98930 51706
rect 98982 51654 98994 51706
rect 99046 51654 99058 51706
rect 99110 51654 99122 51706
rect 99174 51654 99186 51706
rect 99238 51654 100832 51706
rect 97980 51632 100832 51654
rect 1104 51162 1932 51184
rect 1104 51110 1690 51162
rect 1742 51110 1754 51162
rect 1806 51110 1932 51162
rect 1104 51088 1932 51110
rect 97980 51162 100832 51184
rect 97980 51110 99666 51162
rect 99718 51110 99730 51162
rect 99782 51110 99794 51162
rect 99846 51110 99858 51162
rect 99910 51110 99922 51162
rect 99974 51110 100832 51162
rect 97980 51088 100832 51110
rect 1104 50618 1932 50640
rect 1104 50566 1322 50618
rect 1374 50566 1386 50618
rect 1438 50566 1932 50618
rect 1104 50544 1932 50566
rect 97980 50618 100832 50640
rect 97980 50566 98930 50618
rect 98982 50566 98994 50618
rect 99046 50566 99058 50618
rect 99110 50566 99122 50618
rect 99174 50566 99186 50618
rect 99238 50566 100832 50618
rect 97980 50544 100832 50566
rect 1104 50074 1932 50096
rect 1104 50022 1690 50074
rect 1742 50022 1754 50074
rect 1806 50022 1932 50074
rect 1104 50000 1932 50022
rect 97980 50074 100832 50096
rect 97980 50022 99666 50074
rect 99718 50022 99730 50074
rect 99782 50022 99794 50074
rect 99846 50022 99858 50074
rect 99910 50022 99922 50074
rect 99974 50022 100832 50074
rect 97980 50000 100832 50022
rect 1104 49530 1932 49552
rect 1104 49478 1322 49530
rect 1374 49478 1386 49530
rect 1438 49478 1932 49530
rect 1104 49456 1932 49478
rect 97980 49530 100832 49552
rect 97980 49478 98930 49530
rect 98982 49478 98994 49530
rect 99046 49478 99058 49530
rect 99110 49478 99122 49530
rect 99174 49478 99186 49530
rect 99238 49478 100832 49530
rect 97980 49456 100832 49478
rect 1104 48986 1932 49008
rect 1104 48934 1690 48986
rect 1742 48934 1754 48986
rect 1806 48934 1932 48986
rect 1104 48912 1932 48934
rect 97980 48986 100832 49008
rect 97980 48934 99666 48986
rect 99718 48934 99730 48986
rect 99782 48934 99794 48986
rect 99846 48934 99858 48986
rect 99910 48934 99922 48986
rect 99974 48934 100832 48986
rect 97980 48912 100832 48934
rect 1104 48442 1932 48464
rect 1104 48390 1322 48442
rect 1374 48390 1386 48442
rect 1438 48390 1932 48442
rect 1104 48368 1932 48390
rect 97980 48442 100832 48464
rect 97980 48390 98930 48442
rect 98982 48390 98994 48442
rect 99046 48390 99058 48442
rect 99110 48390 99122 48442
rect 99174 48390 99186 48442
rect 99238 48390 100832 48442
rect 97980 48368 100832 48390
rect 1104 47898 1932 47920
rect 1104 47846 1690 47898
rect 1742 47846 1754 47898
rect 1806 47846 1932 47898
rect 1104 47824 1932 47846
rect 97980 47898 100832 47920
rect 97980 47846 99666 47898
rect 99718 47846 99730 47898
rect 99782 47846 99794 47898
rect 99846 47846 99858 47898
rect 99910 47846 99922 47898
rect 99974 47846 100832 47898
rect 97980 47824 100832 47846
rect 1104 47354 1932 47376
rect 1104 47302 1322 47354
rect 1374 47302 1386 47354
rect 1438 47302 1932 47354
rect 1104 47280 1932 47302
rect 97980 47354 100832 47376
rect 97980 47302 98930 47354
rect 98982 47302 98994 47354
rect 99046 47302 99058 47354
rect 99110 47302 99122 47354
rect 99174 47302 99186 47354
rect 99238 47302 100832 47354
rect 97980 47280 100832 47302
rect 1104 46810 1932 46832
rect 1104 46758 1690 46810
rect 1742 46758 1754 46810
rect 1806 46758 1932 46810
rect 1104 46736 1932 46758
rect 97980 46810 100832 46832
rect 97980 46758 99666 46810
rect 99718 46758 99730 46810
rect 99782 46758 99794 46810
rect 99846 46758 99858 46810
rect 99910 46758 99922 46810
rect 99974 46758 100832 46810
rect 97980 46736 100832 46758
rect 1104 46266 1932 46288
rect 1104 46214 1322 46266
rect 1374 46214 1386 46266
rect 1438 46214 1932 46266
rect 1104 46192 1932 46214
rect 97980 46266 100832 46288
rect 97980 46214 98930 46266
rect 98982 46214 98994 46266
rect 99046 46214 99058 46266
rect 99110 46214 99122 46266
rect 99174 46214 99186 46266
rect 99238 46214 100832 46266
rect 97980 46192 100832 46214
rect 98546 46044 98552 46096
rect 98604 46044 98610 46096
rect 98270 45908 98276 45960
rect 98328 45908 98334 45960
rect 98362 45908 98368 45960
rect 98420 45908 98426 45960
rect 98178 45840 98184 45892
rect 98236 45880 98242 45892
rect 98549 45883 98607 45889
rect 98549 45880 98561 45883
rect 98236 45852 98561 45880
rect 98236 45840 98242 45852
rect 98549 45849 98561 45852
rect 98595 45849 98607 45883
rect 98549 45843 98607 45849
rect 1104 45722 1932 45744
rect 1104 45670 1690 45722
rect 1742 45670 1754 45722
rect 1806 45670 1932 45722
rect 1104 45648 1932 45670
rect 97980 45722 100832 45744
rect 97980 45670 99666 45722
rect 99718 45670 99730 45722
rect 99782 45670 99794 45722
rect 99846 45670 99858 45722
rect 99910 45670 99922 45722
rect 99974 45670 100832 45722
rect 97980 45648 100832 45670
rect 1104 45178 1932 45200
rect 1104 45126 1322 45178
rect 1374 45126 1386 45178
rect 1438 45126 1932 45178
rect 1104 45104 1932 45126
rect 97980 45178 100832 45200
rect 97980 45126 98930 45178
rect 98982 45126 98994 45178
rect 99046 45126 99058 45178
rect 99110 45126 99122 45178
rect 99174 45126 99186 45178
rect 99238 45126 100832 45178
rect 97980 45104 100832 45126
rect 98270 45024 98276 45076
rect 98328 45064 98334 45076
rect 98457 45067 98515 45073
rect 98457 45064 98469 45067
rect 98328 45036 98469 45064
rect 98328 45024 98334 45036
rect 98457 45033 98469 45036
rect 98503 45033 98515 45067
rect 98457 45027 98515 45033
rect 98273 44795 98331 44801
rect 98273 44761 98285 44795
rect 98319 44792 98331 44795
rect 98362 44792 98368 44804
rect 98319 44764 98368 44792
rect 98319 44761 98331 44764
rect 98273 44755 98331 44761
rect 98362 44752 98368 44764
rect 98420 44752 98426 44804
rect 98178 44684 98184 44736
rect 98236 44724 98242 44736
rect 98457 44727 98515 44733
rect 98457 44724 98469 44727
rect 98236 44696 98469 44724
rect 98236 44684 98242 44696
rect 98457 44693 98469 44696
rect 98503 44693 98515 44727
rect 98457 44687 98515 44693
rect 98638 44684 98644 44736
rect 98696 44684 98702 44736
rect 1104 44634 1932 44656
rect 1104 44582 1690 44634
rect 1742 44582 1754 44634
rect 1806 44582 1932 44634
rect 1104 44560 1932 44582
rect 97980 44634 100832 44656
rect 97980 44582 99666 44634
rect 99718 44582 99730 44634
rect 99782 44582 99794 44634
rect 99846 44582 99858 44634
rect 99910 44582 99922 44634
rect 99974 44582 100832 44634
rect 97980 44560 100832 44582
rect 1104 44090 1932 44112
rect 1104 44038 1322 44090
rect 1374 44038 1386 44090
rect 1438 44038 1932 44090
rect 1104 44016 1932 44038
rect 97980 44090 100832 44112
rect 97980 44038 98930 44090
rect 98982 44038 98994 44090
rect 99046 44038 99058 44090
rect 99110 44038 99122 44090
rect 99174 44038 99186 44090
rect 99238 44038 100832 44090
rect 97980 44016 100832 44038
rect 1104 43546 1932 43568
rect 1104 43494 1690 43546
rect 1742 43494 1754 43546
rect 1806 43494 1932 43546
rect 1104 43472 1932 43494
rect 97980 43546 100832 43568
rect 97980 43494 99666 43546
rect 99718 43494 99730 43546
rect 99782 43494 99794 43546
rect 99846 43494 99858 43546
rect 99910 43494 99922 43546
rect 99974 43494 100832 43546
rect 97980 43472 100832 43494
rect 97442 43256 97448 43308
rect 97500 43296 97506 43308
rect 98270 43296 98276 43308
rect 97500 43268 98276 43296
rect 97500 43256 97506 43268
rect 98270 43256 98276 43268
rect 98328 43256 98334 43308
rect 98362 43052 98368 43104
rect 98420 43052 98426 43104
rect 1104 43002 1932 43024
rect 1104 42950 1322 43002
rect 1374 42950 1386 43002
rect 1438 42950 1932 43002
rect 1104 42928 1932 42950
rect 97980 43002 100832 43024
rect 97980 42950 98930 43002
rect 98982 42950 98994 43002
rect 99046 42950 99058 43002
rect 99110 42950 99122 43002
rect 99174 42950 99186 43002
rect 99238 42950 100832 43002
rect 97980 42928 100832 42950
rect 1104 42458 1932 42480
rect 1104 42406 1690 42458
rect 1742 42406 1754 42458
rect 1806 42406 1932 42458
rect 1104 42384 1932 42406
rect 97980 42458 100832 42480
rect 97980 42406 99666 42458
rect 99718 42406 99730 42458
rect 99782 42406 99794 42458
rect 99846 42406 99858 42458
rect 99910 42406 99922 42458
rect 99974 42406 100832 42458
rect 97980 42384 100832 42406
rect 1104 41914 1932 41936
rect 1104 41862 1322 41914
rect 1374 41862 1386 41914
rect 1438 41862 1932 41914
rect 1104 41840 1932 41862
rect 97980 41914 100832 41936
rect 97980 41862 98930 41914
rect 98982 41862 98994 41914
rect 99046 41862 99058 41914
rect 99110 41862 99122 41914
rect 99174 41862 99186 41914
rect 99238 41862 100832 41914
rect 97980 41840 100832 41862
rect 1104 41370 1932 41392
rect 1104 41318 1690 41370
rect 1742 41318 1754 41370
rect 1806 41318 1932 41370
rect 1104 41296 1932 41318
rect 97980 41370 100832 41392
rect 97980 41318 99666 41370
rect 99718 41318 99730 41370
rect 99782 41318 99794 41370
rect 99846 41318 99858 41370
rect 99910 41318 99922 41370
rect 99974 41318 100832 41370
rect 97980 41296 100832 41318
rect 98362 41148 98368 41200
rect 98420 41188 98426 41200
rect 98420 41160 98670 41188
rect 98420 41148 98426 41160
rect 98454 41012 98460 41064
rect 98512 41052 98518 41064
rect 99837 41055 99895 41061
rect 99837 41052 99849 41055
rect 98512 41024 99849 41052
rect 98512 41012 98518 41024
rect 99837 41021 99849 41024
rect 99883 41021 99895 41055
rect 99837 41015 99895 41021
rect 100110 41012 100116 41064
rect 100168 41012 100174 41064
rect 98178 40876 98184 40928
rect 98236 40916 98242 40928
rect 98365 40919 98423 40925
rect 98365 40916 98377 40919
rect 98236 40888 98377 40916
rect 98236 40876 98242 40888
rect 98365 40885 98377 40888
rect 98411 40885 98423 40919
rect 98365 40879 98423 40885
rect 1104 40826 1932 40848
rect 1104 40774 1322 40826
rect 1374 40774 1386 40826
rect 1438 40774 1932 40826
rect 1104 40752 1932 40774
rect 97980 40826 100832 40848
rect 97980 40774 98930 40826
rect 98982 40774 98994 40826
rect 99046 40774 99058 40826
rect 99110 40774 99122 40826
rect 99174 40774 99186 40826
rect 99238 40774 100832 40826
rect 97980 40752 100832 40774
rect 98454 40672 98460 40724
rect 98512 40672 98518 40724
rect 98273 40511 98331 40517
rect 98273 40477 98285 40511
rect 98319 40477 98331 40511
rect 98273 40471 98331 40477
rect 98457 40511 98515 40517
rect 98457 40477 98469 40511
rect 98503 40508 98515 40511
rect 98546 40508 98552 40520
rect 98503 40480 98552 40508
rect 98503 40477 98515 40480
rect 98457 40471 98515 40477
rect 98288 40440 98316 40471
rect 98546 40468 98552 40480
rect 98604 40468 98610 40520
rect 98638 40440 98644 40452
rect 98288 40412 98644 40440
rect 98638 40400 98644 40412
rect 98696 40440 98702 40452
rect 100202 40440 100208 40452
rect 98696 40412 100208 40440
rect 98696 40400 98702 40412
rect 100202 40400 100208 40412
rect 100260 40400 100266 40452
rect 1104 40282 1932 40304
rect 1104 40230 1690 40282
rect 1742 40230 1754 40282
rect 1806 40230 1932 40282
rect 1104 40208 1932 40230
rect 97980 40282 100832 40304
rect 97980 40230 99666 40282
rect 99718 40230 99730 40282
rect 99782 40230 99794 40282
rect 99846 40230 99858 40282
rect 99910 40230 99922 40282
rect 99974 40230 100832 40282
rect 97980 40208 100832 40230
rect 1104 39738 1932 39760
rect 1104 39686 1322 39738
rect 1374 39686 1386 39738
rect 1438 39686 1932 39738
rect 1104 39664 1932 39686
rect 97980 39738 100832 39760
rect 97980 39686 98930 39738
rect 98982 39686 98994 39738
rect 99046 39686 99058 39738
rect 99110 39686 99122 39738
rect 99174 39686 99186 39738
rect 99238 39686 100832 39738
rect 97980 39664 100832 39686
rect 1104 39194 1932 39216
rect 1104 39142 1690 39194
rect 1742 39142 1754 39194
rect 1806 39142 1932 39194
rect 1104 39120 1932 39142
rect 97980 39194 100832 39216
rect 97980 39142 99666 39194
rect 99718 39142 99730 39194
rect 99782 39142 99794 39194
rect 99846 39142 99858 39194
rect 99910 39142 99922 39194
rect 99974 39142 100832 39194
rect 97980 39120 100832 39142
rect 1104 38650 1932 38672
rect 1104 38598 1322 38650
rect 1374 38598 1386 38650
rect 1438 38598 1932 38650
rect 1104 38576 1932 38598
rect 97980 38650 100832 38672
rect 97980 38598 98930 38650
rect 98982 38598 98994 38650
rect 99046 38598 99058 38650
rect 99110 38598 99122 38650
rect 99174 38598 99186 38650
rect 99238 38598 100832 38650
rect 97980 38576 100832 38598
rect 1104 38106 1932 38128
rect 1104 38054 1690 38106
rect 1742 38054 1754 38106
rect 1806 38054 1932 38106
rect 1104 38032 1932 38054
rect 97980 38106 100832 38128
rect 97980 38054 99666 38106
rect 99718 38054 99730 38106
rect 99782 38054 99794 38106
rect 99846 38054 99858 38106
rect 99910 38054 99922 38106
rect 99974 38054 100832 38106
rect 97980 38032 100832 38054
rect 1104 37562 1932 37584
rect 1104 37510 1322 37562
rect 1374 37510 1386 37562
rect 1438 37510 1932 37562
rect 1104 37488 1932 37510
rect 97980 37562 100832 37584
rect 97980 37510 98930 37562
rect 98982 37510 98994 37562
rect 99046 37510 99058 37562
rect 99110 37510 99122 37562
rect 99174 37510 99186 37562
rect 99238 37510 100832 37562
rect 97980 37488 100832 37510
rect 1104 37018 1932 37040
rect 1104 36966 1690 37018
rect 1742 36966 1754 37018
rect 1806 36966 1932 37018
rect 1104 36944 1932 36966
rect 97980 37018 100832 37040
rect 97980 36966 99666 37018
rect 99718 36966 99730 37018
rect 99782 36966 99794 37018
rect 99846 36966 99858 37018
rect 99910 36966 99922 37018
rect 99974 36966 100832 37018
rect 97980 36944 100832 36966
rect 1104 36474 1932 36496
rect 1104 36422 1322 36474
rect 1374 36422 1386 36474
rect 1438 36422 1932 36474
rect 1104 36400 1932 36422
rect 97980 36474 100832 36496
rect 97980 36422 98930 36474
rect 98982 36422 98994 36474
rect 99046 36422 99058 36474
rect 99110 36422 99122 36474
rect 99174 36422 99186 36474
rect 99238 36422 100832 36474
rect 97980 36400 100832 36422
rect 1104 35930 1932 35952
rect 1104 35878 1690 35930
rect 1742 35878 1754 35930
rect 1806 35878 1932 35930
rect 1104 35856 1932 35878
rect 97980 35930 100832 35952
rect 97980 35878 99666 35930
rect 99718 35878 99730 35930
rect 99782 35878 99794 35930
rect 99846 35878 99858 35930
rect 99910 35878 99922 35930
rect 99974 35878 100832 35930
rect 97980 35856 100832 35878
rect 98270 35640 98276 35692
rect 98328 35680 98334 35692
rect 98454 35680 98460 35692
rect 98328 35652 98460 35680
rect 98328 35640 98334 35652
rect 98454 35640 98460 35652
rect 98512 35640 98518 35692
rect 98365 35479 98423 35485
rect 98365 35445 98377 35479
rect 98411 35476 98423 35479
rect 98730 35476 98736 35488
rect 98411 35448 98736 35476
rect 98411 35445 98423 35448
rect 98365 35439 98423 35445
rect 98730 35436 98736 35448
rect 98788 35436 98794 35488
rect 1104 35386 1932 35408
rect 1104 35334 1322 35386
rect 1374 35334 1386 35386
rect 1438 35334 1932 35386
rect 1104 35312 1932 35334
rect 97980 35386 100832 35408
rect 97980 35334 98930 35386
rect 98982 35334 98994 35386
rect 99046 35334 99058 35386
rect 99110 35334 99122 35386
rect 99174 35334 99186 35386
rect 99238 35334 100832 35386
rect 97980 35312 100832 35334
rect 1104 34842 1932 34864
rect 1104 34790 1690 34842
rect 1742 34790 1754 34842
rect 1806 34790 1932 34842
rect 1104 34768 1932 34790
rect 97980 34842 100832 34864
rect 97980 34790 99666 34842
rect 99718 34790 99730 34842
rect 99782 34790 99794 34842
rect 99846 34790 99858 34842
rect 99910 34790 99922 34842
rect 99974 34790 100832 34842
rect 97980 34768 100832 34790
rect 98273 34595 98331 34601
rect 98273 34561 98285 34595
rect 98319 34592 98331 34595
rect 98454 34592 98460 34604
rect 98319 34564 98460 34592
rect 98319 34561 98331 34564
rect 98273 34555 98331 34561
rect 98454 34552 98460 34564
rect 98512 34552 98518 34604
rect 98362 34484 98368 34536
rect 98420 34484 98426 34536
rect 1104 34298 1932 34320
rect 1104 34246 1322 34298
rect 1374 34246 1386 34298
rect 1438 34246 1932 34298
rect 1104 34224 1932 34246
rect 97980 34298 100832 34320
rect 97980 34246 98930 34298
rect 98982 34246 98994 34298
rect 99046 34246 99058 34298
rect 99110 34246 99122 34298
rect 99174 34246 99186 34298
rect 99238 34246 100832 34298
rect 97980 34224 100832 34246
rect 1104 33754 1932 33776
rect 1104 33702 1690 33754
rect 1742 33702 1754 33754
rect 1806 33702 1932 33754
rect 1104 33680 1932 33702
rect 97980 33754 100832 33776
rect 97980 33702 99666 33754
rect 99718 33702 99730 33754
rect 99782 33702 99794 33754
rect 99846 33702 99858 33754
rect 99910 33702 99922 33754
rect 99974 33702 100832 33754
rect 97980 33680 100832 33702
rect 1104 33210 1932 33232
rect 1104 33158 1322 33210
rect 1374 33158 1386 33210
rect 1438 33158 1932 33210
rect 1104 33136 1932 33158
rect 97980 33210 100832 33232
rect 97980 33158 98930 33210
rect 98982 33158 98994 33210
rect 99046 33158 99058 33210
rect 99110 33158 99122 33210
rect 99174 33158 99186 33210
rect 99238 33158 100832 33210
rect 97980 33136 100832 33158
rect 1104 32666 1932 32688
rect 1104 32614 1690 32666
rect 1742 32614 1754 32666
rect 1806 32614 1932 32666
rect 1104 32592 1932 32614
rect 97980 32666 100832 32688
rect 97980 32614 99666 32666
rect 99718 32614 99730 32666
rect 99782 32614 99794 32666
rect 99846 32614 99858 32666
rect 99910 32614 99922 32666
rect 99974 32614 100832 32666
rect 97980 32592 100832 32614
rect 1104 32122 1932 32144
rect 1104 32070 1322 32122
rect 1374 32070 1386 32122
rect 1438 32070 1932 32122
rect 1104 32048 1932 32070
rect 97980 32122 100832 32144
rect 97980 32070 98930 32122
rect 98982 32070 98994 32122
rect 99046 32070 99058 32122
rect 99110 32070 99122 32122
rect 99174 32070 99186 32122
rect 99238 32070 100832 32122
rect 97980 32048 100832 32070
rect 98365 31875 98423 31881
rect 98365 31841 98377 31875
rect 98411 31872 98423 31875
rect 99374 31872 99380 31884
rect 98411 31844 99380 31872
rect 98411 31841 98423 31844
rect 98365 31835 98423 31841
rect 99374 31832 99380 31844
rect 99432 31832 99438 31884
rect 99834 31832 99840 31884
rect 99892 31832 99898 31884
rect 98730 31764 98736 31816
rect 98788 31764 98794 31816
rect 100113 31807 100171 31813
rect 100113 31773 100125 31807
rect 100159 31804 100171 31807
rect 100202 31804 100208 31816
rect 100159 31776 100208 31804
rect 100159 31773 100171 31776
rect 100113 31767 100171 31773
rect 100202 31764 100208 31776
rect 100260 31764 100266 31816
rect 1104 31578 1932 31600
rect 1104 31526 1690 31578
rect 1742 31526 1754 31578
rect 1806 31526 1932 31578
rect 1104 31504 1932 31526
rect 97980 31578 100832 31600
rect 97980 31526 99666 31578
rect 99718 31526 99730 31578
rect 99782 31526 99794 31578
rect 99846 31526 99858 31578
rect 99910 31526 99922 31578
rect 99974 31526 100832 31578
rect 97980 31504 100832 31526
rect 1104 31034 1932 31056
rect 1104 30982 1322 31034
rect 1374 30982 1386 31034
rect 1438 30982 1932 31034
rect 1104 30960 1932 30982
rect 97980 31034 100832 31056
rect 97980 30982 98930 31034
rect 98982 30982 98994 31034
rect 99046 30982 99058 31034
rect 99110 30982 99122 31034
rect 99174 30982 99186 31034
rect 99238 30982 100832 31034
rect 97980 30960 100832 30982
rect 100021 30719 100079 30725
rect 100021 30685 100033 30719
rect 100067 30716 100079 30719
rect 100202 30716 100208 30728
rect 100067 30688 100208 30716
rect 100067 30685 100079 30688
rect 100021 30679 100079 30685
rect 100202 30676 100208 30688
rect 100260 30676 100266 30728
rect 98362 30608 98368 30660
rect 98420 30648 98426 30660
rect 99745 30651 99803 30657
rect 98420 30620 98578 30648
rect 98420 30608 98426 30620
rect 99745 30617 99757 30651
rect 99791 30617 99803 30651
rect 99745 30611 99803 30617
rect 98270 30540 98276 30592
rect 98328 30540 98334 30592
rect 99558 30540 99564 30592
rect 99616 30580 99622 30592
rect 99760 30580 99788 30611
rect 99616 30552 99788 30580
rect 99616 30540 99622 30552
rect 1104 30490 1932 30512
rect 1104 30438 1690 30490
rect 1742 30438 1754 30490
rect 1806 30438 1932 30490
rect 1104 30416 1932 30438
rect 97980 30490 100832 30512
rect 97980 30438 99666 30490
rect 99718 30438 99730 30490
rect 99782 30438 99794 30490
rect 99846 30438 99858 30490
rect 99910 30438 99922 30490
rect 99974 30438 100832 30490
rect 97980 30416 100832 30438
rect 98825 30243 98883 30249
rect 98825 30209 98837 30243
rect 98871 30240 98883 30243
rect 99374 30240 99380 30252
rect 98871 30212 99380 30240
rect 98871 30209 98883 30212
rect 98825 30203 98883 30209
rect 99374 30200 99380 30212
rect 99432 30240 99438 30252
rect 100110 30240 100116 30252
rect 99432 30212 100116 30240
rect 99432 30200 99438 30212
rect 100110 30200 100116 30212
rect 100168 30200 100174 30252
rect 99374 29996 99380 30048
rect 99432 29996 99438 30048
rect 1104 29946 1932 29968
rect 1104 29894 1322 29946
rect 1374 29894 1386 29946
rect 1438 29894 1932 29946
rect 1104 29872 1932 29894
rect 97980 29946 100832 29968
rect 97980 29894 98930 29946
rect 98982 29894 98994 29946
rect 99046 29894 99058 29946
rect 99110 29894 99122 29946
rect 99174 29894 99186 29946
rect 99238 29894 100832 29946
rect 97980 29872 100832 29894
rect 98273 29631 98331 29637
rect 98273 29597 98285 29631
rect 98319 29628 98331 29631
rect 98454 29628 98460 29640
rect 98319 29600 98460 29628
rect 98319 29597 98331 29600
rect 98273 29591 98331 29597
rect 98454 29588 98460 29600
rect 98512 29628 98518 29640
rect 98730 29628 98736 29640
rect 98512 29600 98736 29628
rect 98512 29588 98518 29600
rect 98730 29588 98736 29600
rect 98788 29588 98794 29640
rect 98365 29495 98423 29501
rect 98365 29461 98377 29495
rect 98411 29492 98423 29495
rect 98638 29492 98644 29504
rect 98411 29464 98644 29492
rect 98411 29461 98423 29464
rect 98365 29455 98423 29461
rect 98638 29452 98644 29464
rect 98696 29452 98702 29504
rect 1104 29402 1932 29424
rect 1104 29350 1690 29402
rect 1742 29350 1754 29402
rect 1806 29350 1932 29402
rect 1104 29328 1932 29350
rect 97980 29402 100832 29424
rect 97980 29350 99666 29402
rect 99718 29350 99730 29402
rect 99782 29350 99794 29402
rect 99846 29350 99858 29402
rect 99910 29350 99922 29402
rect 99974 29350 100832 29402
rect 97980 29328 100832 29350
rect 98365 29155 98423 29161
rect 98365 29121 98377 29155
rect 98411 29152 98423 29155
rect 98730 29152 98736 29164
rect 98411 29124 98736 29152
rect 98411 29121 98423 29124
rect 98365 29115 98423 29121
rect 98730 29112 98736 29124
rect 98788 29112 98794 29164
rect 99374 29112 99380 29164
rect 99432 29152 99438 29164
rect 99929 29155 99987 29161
rect 99929 29152 99941 29155
rect 99432 29124 99941 29152
rect 99432 29112 99438 29124
rect 99929 29121 99941 29124
rect 99975 29121 99987 29155
rect 99929 29115 99987 29121
rect 98270 29044 98276 29096
rect 98328 29084 98334 29096
rect 98917 29087 98975 29093
rect 98917 29084 98929 29087
rect 98328 29056 98929 29084
rect 98328 29044 98334 29056
rect 98917 29053 98929 29056
rect 98963 29084 98975 29087
rect 99282 29084 99288 29096
rect 98963 29056 99288 29084
rect 98963 29053 98975 29056
rect 98917 29047 98975 29053
rect 99282 29044 99288 29056
rect 99340 29044 99346 29096
rect 99837 29087 99895 29093
rect 99837 29053 99849 29087
rect 99883 29084 99895 29087
rect 100294 29084 100300 29096
rect 99883 29056 100300 29084
rect 99883 29053 99895 29056
rect 99837 29047 99895 29053
rect 100294 29044 100300 29056
rect 100352 29044 100358 29096
rect 98457 29019 98515 29025
rect 98457 28985 98469 29019
rect 98503 29016 98515 29019
rect 98546 29016 98552 29028
rect 98503 28988 98552 29016
rect 98503 28985 98515 28988
rect 98457 28979 98515 28985
rect 98546 28976 98552 28988
rect 98604 28976 98610 29028
rect 99466 28976 99472 29028
rect 99524 28976 99530 29028
rect 99561 29019 99619 29025
rect 99561 28985 99573 29019
rect 99607 29016 99619 29019
rect 100018 29016 100024 29028
rect 99607 28988 100024 29016
rect 99607 28985 99619 28988
rect 99561 28979 99619 28985
rect 100018 28976 100024 28988
rect 100076 28976 100082 29028
rect 1104 28858 1932 28880
rect 1104 28806 1322 28858
rect 1374 28806 1386 28858
rect 1438 28806 1932 28858
rect 1104 28784 1932 28806
rect 97980 28858 100832 28880
rect 97980 28806 98930 28858
rect 98982 28806 98994 28858
rect 99046 28806 99058 28858
rect 99110 28806 99122 28858
rect 99174 28806 99186 28858
rect 99238 28806 100832 28858
rect 97980 28784 100832 28806
rect 1104 28314 1932 28336
rect 1104 28262 1690 28314
rect 1742 28262 1754 28314
rect 1806 28262 1932 28314
rect 1104 28240 1932 28262
rect 97980 28314 100832 28336
rect 97980 28262 99666 28314
rect 99718 28262 99730 28314
rect 99782 28262 99794 28314
rect 99846 28262 99858 28314
rect 99910 28262 99922 28314
rect 99974 28262 100832 28314
rect 97980 28240 100832 28262
rect 1104 27770 1932 27792
rect 1104 27718 1322 27770
rect 1374 27718 1386 27770
rect 1438 27718 1932 27770
rect 1104 27696 1932 27718
rect 97980 27770 100832 27792
rect 97980 27718 98930 27770
rect 98982 27718 98994 27770
rect 99046 27718 99058 27770
rect 99110 27718 99122 27770
rect 99174 27718 99186 27770
rect 99238 27718 100832 27770
rect 97980 27696 100832 27718
rect 97350 27548 97356 27600
rect 97408 27588 97414 27600
rect 98362 27588 98368 27600
rect 97408 27560 98368 27588
rect 97408 27548 97414 27560
rect 98362 27548 98368 27560
rect 98420 27548 98426 27600
rect 99558 27548 99564 27600
rect 99616 27588 99622 27600
rect 99653 27591 99711 27597
rect 99653 27588 99665 27591
rect 99616 27560 99665 27588
rect 99616 27548 99622 27560
rect 99653 27557 99665 27560
rect 99699 27557 99711 27591
rect 99653 27551 99711 27557
rect 99377 27523 99435 27529
rect 99377 27489 99389 27523
rect 99423 27520 99435 27523
rect 99837 27523 99895 27529
rect 99837 27520 99849 27523
rect 99423 27492 99849 27520
rect 99423 27489 99435 27492
rect 99377 27483 99435 27489
rect 99837 27489 99849 27492
rect 99883 27489 99895 27523
rect 99837 27483 99895 27489
rect 99285 27455 99343 27461
rect 99285 27421 99297 27455
rect 99331 27452 99343 27455
rect 99466 27452 99472 27464
rect 99331 27424 99472 27452
rect 99331 27421 99343 27424
rect 99285 27415 99343 27421
rect 99466 27412 99472 27424
rect 99524 27412 99530 27464
rect 99745 27455 99803 27461
rect 99745 27421 99757 27455
rect 99791 27421 99803 27455
rect 99745 27415 99803 27421
rect 99929 27455 99987 27461
rect 99929 27421 99941 27455
rect 99975 27452 99987 27455
rect 100018 27452 100024 27464
rect 99975 27424 100024 27452
rect 99975 27421 99987 27424
rect 99929 27415 99987 27421
rect 99558 27344 99564 27396
rect 99616 27384 99622 27396
rect 99760 27384 99788 27415
rect 100018 27412 100024 27424
rect 100076 27452 100082 27464
rect 100294 27452 100300 27464
rect 100076 27424 100300 27452
rect 100076 27412 100082 27424
rect 100294 27412 100300 27424
rect 100352 27412 100358 27464
rect 100110 27384 100116 27396
rect 99616 27356 100116 27384
rect 99616 27344 99622 27356
rect 100110 27344 100116 27356
rect 100168 27344 100174 27396
rect 1104 27226 1932 27248
rect 1104 27174 1690 27226
rect 1742 27174 1754 27226
rect 1806 27174 1932 27226
rect 1104 27152 1932 27174
rect 97980 27226 100832 27248
rect 97980 27174 99666 27226
rect 99718 27174 99730 27226
rect 99782 27174 99794 27226
rect 99846 27174 99858 27226
rect 99910 27174 99922 27226
rect 99974 27174 100832 27226
rect 97980 27152 100832 27174
rect 1104 26682 1932 26704
rect 1104 26630 1322 26682
rect 1374 26630 1386 26682
rect 1438 26630 1932 26682
rect 1104 26608 1932 26630
rect 97980 26682 100832 26704
rect 97980 26630 98930 26682
rect 98982 26630 98994 26682
rect 99046 26630 99058 26682
rect 99110 26630 99122 26682
rect 99174 26630 99186 26682
rect 99238 26630 100832 26682
rect 97980 26608 100832 26630
rect 100297 26503 100355 26509
rect 100297 26469 100309 26503
rect 100343 26469 100355 26503
rect 100297 26463 100355 26469
rect 98362 26392 98368 26444
rect 98420 26432 98426 26444
rect 98641 26435 98699 26441
rect 98641 26432 98653 26435
rect 98420 26404 98653 26432
rect 98420 26392 98426 26404
rect 98641 26401 98653 26404
rect 98687 26401 98699 26435
rect 98641 26395 98699 26401
rect 98917 26367 98975 26373
rect 98917 26333 98929 26367
rect 98963 26364 98975 26367
rect 100312 26364 100340 26463
rect 98963 26336 100340 26364
rect 98963 26333 98975 26336
rect 98917 26327 98975 26333
rect 100478 26324 100484 26376
rect 100536 26324 100542 26376
rect 1104 26138 1932 26160
rect 1104 26086 1690 26138
rect 1742 26086 1754 26138
rect 1806 26086 1932 26138
rect 1104 26064 1932 26086
rect 97980 26138 100832 26160
rect 97980 26086 99666 26138
rect 99718 26086 99730 26138
rect 99782 26086 99794 26138
rect 99846 26086 99858 26138
rect 99910 26086 99922 26138
rect 99974 26086 100832 26138
rect 97980 26064 100832 26086
rect 99540 26027 99598 26033
rect 99540 25993 99552 26027
rect 99586 26024 99598 26027
rect 100018 26024 100024 26036
rect 99586 25996 100024 26024
rect 99586 25993 99598 25996
rect 99540 25987 99598 25993
rect 100018 25984 100024 25996
rect 100076 25984 100082 26036
rect 98362 25916 98368 25968
rect 98420 25916 98426 25968
rect 99745 25959 99803 25965
rect 99745 25956 99757 25959
rect 99576 25928 99757 25956
rect 99576 25900 99604 25928
rect 99745 25925 99757 25928
rect 99791 25925 99803 25959
rect 99745 25919 99803 25925
rect 99558 25848 99564 25900
rect 99616 25848 99622 25900
rect 98362 25780 98368 25832
rect 98420 25820 98426 25832
rect 98730 25820 98736 25832
rect 98420 25792 98736 25820
rect 98420 25780 98426 25792
rect 98730 25780 98736 25792
rect 98788 25820 98794 25832
rect 99101 25823 99159 25829
rect 99101 25820 99113 25823
rect 98788 25792 99113 25820
rect 98788 25780 98794 25792
rect 99101 25789 99113 25792
rect 99147 25789 99159 25823
rect 99101 25783 99159 25789
rect 98822 25712 98828 25764
rect 98880 25752 98886 25764
rect 99282 25752 99288 25764
rect 98880 25724 99288 25752
rect 98880 25712 98886 25724
rect 99282 25712 99288 25724
rect 99340 25752 99346 25764
rect 99340 25724 99604 25752
rect 99340 25712 99346 25724
rect 98270 25644 98276 25696
rect 98328 25684 98334 25696
rect 99576 25693 99604 25724
rect 99377 25687 99435 25693
rect 99377 25684 99389 25687
rect 98328 25656 99389 25684
rect 98328 25644 98334 25656
rect 99377 25653 99389 25656
rect 99423 25653 99435 25687
rect 99377 25647 99435 25653
rect 99561 25687 99619 25693
rect 99561 25653 99573 25687
rect 99607 25653 99619 25687
rect 99561 25647 99619 25653
rect 1104 25594 1932 25616
rect 1104 25542 1322 25594
rect 1374 25542 1386 25594
rect 1438 25542 1932 25594
rect 1104 25520 1932 25542
rect 97980 25594 100832 25616
rect 97980 25542 98930 25594
rect 98982 25542 98994 25594
rect 99046 25542 99058 25594
rect 99110 25542 99122 25594
rect 99174 25542 99186 25594
rect 99238 25542 100832 25594
rect 97980 25520 100832 25542
rect 98638 25304 98644 25356
rect 98696 25304 98702 25356
rect 99282 25304 99288 25356
rect 99340 25344 99346 25356
rect 99837 25347 99895 25353
rect 99837 25344 99849 25347
rect 99340 25316 99849 25344
rect 99340 25304 99346 25316
rect 99837 25313 99849 25316
rect 99883 25313 99895 25347
rect 99837 25307 99895 25313
rect 98656 25276 98684 25304
rect 100113 25279 100171 25285
rect 98656 25248 98762 25276
rect 100113 25245 100125 25279
rect 100159 25276 100171 25279
rect 100202 25276 100208 25288
rect 100159 25248 100208 25276
rect 100159 25245 100171 25248
rect 100113 25239 100171 25245
rect 100202 25236 100208 25248
rect 100260 25236 100266 25288
rect 98086 25100 98092 25152
rect 98144 25140 98150 25152
rect 98365 25143 98423 25149
rect 98365 25140 98377 25143
rect 98144 25112 98377 25140
rect 98144 25100 98150 25112
rect 98365 25109 98377 25112
rect 98411 25109 98423 25143
rect 98365 25103 98423 25109
rect 1104 25050 1932 25072
rect 1104 24998 1690 25050
rect 1742 24998 1754 25050
rect 1806 24998 1932 25050
rect 1104 24976 1932 24998
rect 97980 25050 100832 25072
rect 97980 24998 99666 25050
rect 99718 24998 99730 25050
rect 99782 24998 99794 25050
rect 99846 24998 99858 25050
rect 99910 24998 99922 25050
rect 99974 24998 100832 25050
rect 97980 24976 100832 24998
rect 98546 24760 98552 24812
rect 98604 24800 98610 24812
rect 98604 24772 98854 24800
rect 98604 24760 98610 24772
rect 99374 24692 99380 24744
rect 99432 24732 99438 24744
rect 99929 24735 99987 24741
rect 99929 24732 99941 24735
rect 99432 24704 99941 24732
rect 99432 24692 99438 24704
rect 99929 24701 99941 24704
rect 99975 24701 99987 24735
rect 99929 24695 99987 24701
rect 100202 24692 100208 24744
rect 100260 24692 100266 24744
rect 98457 24599 98515 24605
rect 98457 24565 98469 24599
rect 98503 24596 98515 24599
rect 98546 24596 98552 24608
rect 98503 24568 98552 24596
rect 98503 24565 98515 24568
rect 98457 24559 98515 24565
rect 98546 24556 98552 24568
rect 98604 24556 98610 24608
rect 1104 24506 1932 24528
rect 1104 24454 1322 24506
rect 1374 24454 1386 24506
rect 1438 24454 1932 24506
rect 1104 24432 1932 24454
rect 97980 24506 100832 24528
rect 97980 24454 98930 24506
rect 98982 24454 98994 24506
rect 99046 24454 99058 24506
rect 99110 24454 99122 24506
rect 99174 24454 99186 24506
rect 99238 24454 100832 24506
rect 97980 24432 100832 24454
rect 98362 24148 98368 24200
rect 98420 24148 98426 24200
rect 98454 24012 98460 24064
rect 98512 24012 98518 24064
rect 1104 23962 1932 23984
rect 1104 23910 1690 23962
rect 1742 23910 1754 23962
rect 1806 23910 1932 23962
rect 1104 23888 1932 23910
rect 97980 23962 100832 23984
rect 97980 23910 99666 23962
rect 99718 23910 99730 23962
rect 99782 23910 99794 23962
rect 99846 23910 99858 23962
rect 99910 23910 99922 23962
rect 99974 23910 100832 23962
rect 97980 23888 100832 23910
rect 98730 23808 98736 23860
rect 98788 23808 98794 23860
rect 98917 23851 98975 23857
rect 98917 23817 98929 23851
rect 98963 23848 98975 23851
rect 99282 23848 99288 23860
rect 98963 23820 99288 23848
rect 98963 23817 98975 23820
rect 98917 23811 98975 23817
rect 99282 23808 99288 23820
rect 99340 23808 99346 23860
rect 98270 23672 98276 23724
rect 98328 23672 98334 23724
rect 98792 23715 98850 23721
rect 98792 23681 98804 23715
rect 98838 23712 98850 23715
rect 99466 23712 99472 23724
rect 98838 23684 99472 23712
rect 98838 23681 98850 23684
rect 98792 23675 98850 23681
rect 99466 23672 99472 23684
rect 99524 23712 99530 23724
rect 100018 23712 100024 23724
rect 99524 23684 100024 23712
rect 99524 23672 99530 23684
rect 100018 23672 100024 23684
rect 100076 23672 100082 23724
rect 98086 23468 98092 23520
rect 98144 23508 98150 23520
rect 98362 23508 98368 23520
rect 98144 23480 98368 23508
rect 98144 23468 98150 23480
rect 98362 23468 98368 23480
rect 98420 23468 98426 23520
rect 1104 23418 1932 23440
rect 1104 23366 1322 23418
rect 1374 23366 1386 23418
rect 1438 23366 1932 23418
rect 1104 23344 1932 23366
rect 97980 23418 100832 23440
rect 97980 23366 98930 23418
rect 98982 23366 98994 23418
rect 99046 23366 99058 23418
rect 99110 23366 99122 23418
rect 99174 23366 99186 23418
rect 99238 23366 100832 23418
rect 97980 23344 100832 23366
rect 1104 22874 1932 22896
rect 1104 22822 1690 22874
rect 1742 22822 1754 22874
rect 1806 22822 1932 22874
rect 1104 22800 1932 22822
rect 97980 22874 100832 22896
rect 97980 22822 99666 22874
rect 99718 22822 99730 22874
rect 99782 22822 99794 22874
rect 99846 22822 99858 22874
rect 99910 22822 99922 22874
rect 99974 22822 100832 22874
rect 97980 22800 100832 22822
rect 97350 22720 97356 22772
rect 97408 22760 97414 22772
rect 98362 22760 98368 22772
rect 97408 22732 98368 22760
rect 97408 22720 97414 22732
rect 98362 22720 98368 22732
rect 98420 22760 98426 22772
rect 98473 22763 98531 22769
rect 98473 22760 98485 22763
rect 98420 22732 98485 22760
rect 98420 22720 98426 22732
rect 98473 22729 98485 22732
rect 98519 22729 98531 22763
rect 98473 22723 98531 22729
rect 98641 22763 98699 22769
rect 98641 22729 98653 22763
rect 98687 22760 98699 22763
rect 98730 22760 98736 22772
rect 98687 22732 98736 22760
rect 98687 22729 98699 22732
rect 98641 22723 98699 22729
rect 98730 22720 98736 22732
rect 98788 22720 98794 22772
rect 99374 22720 99380 22772
rect 99432 22720 99438 22772
rect 99466 22720 99472 22772
rect 99524 22720 99530 22772
rect 98273 22695 98331 22701
rect 98273 22692 98285 22695
rect 98196 22664 98285 22692
rect 98196 22488 98224 22664
rect 98273 22661 98285 22664
rect 98319 22661 98331 22695
rect 98273 22655 98331 22661
rect 98748 22633 98776 22720
rect 98825 22695 98883 22701
rect 98825 22661 98837 22695
rect 98871 22692 98883 22695
rect 99484 22692 99512 22720
rect 98871 22664 99512 22692
rect 98871 22661 98883 22664
rect 98825 22655 98883 22661
rect 98733 22627 98791 22633
rect 98733 22593 98745 22627
rect 98779 22593 98791 22627
rect 99009 22627 99067 22633
rect 99009 22624 99021 22627
rect 98733 22587 98791 22593
rect 98932 22596 99021 22624
rect 98270 22516 98276 22568
rect 98328 22556 98334 22568
rect 98546 22556 98552 22568
rect 98328 22528 98552 22556
rect 98328 22516 98334 22528
rect 98546 22516 98552 22528
rect 98604 22556 98610 22568
rect 98932 22556 98960 22596
rect 99009 22593 99021 22596
rect 99055 22593 99067 22627
rect 99009 22587 99067 22593
rect 99282 22584 99288 22636
rect 99340 22584 99346 22636
rect 99469 22627 99527 22633
rect 99469 22593 99481 22627
rect 99515 22593 99527 22627
rect 99469 22587 99527 22593
rect 99484 22556 99512 22587
rect 98604 22528 98960 22556
rect 99024 22528 99512 22556
rect 98604 22516 98610 22528
rect 99024 22497 99052 22528
rect 99009 22491 99067 22497
rect 98196 22460 98960 22488
rect 98457 22423 98515 22429
rect 98457 22389 98469 22423
rect 98503 22420 98515 22423
rect 98546 22420 98552 22432
rect 98503 22392 98552 22420
rect 98503 22389 98515 22392
rect 98457 22383 98515 22389
rect 98546 22380 98552 22392
rect 98604 22420 98610 22432
rect 98822 22420 98828 22432
rect 98604 22392 98828 22420
rect 98604 22380 98610 22392
rect 98822 22380 98828 22392
rect 98880 22380 98886 22432
rect 98932 22420 98960 22460
rect 99009 22457 99021 22491
rect 99055 22457 99067 22491
rect 99009 22451 99067 22457
rect 99374 22420 99380 22432
rect 98932 22392 99380 22420
rect 99374 22380 99380 22392
rect 99432 22420 99438 22432
rect 99558 22420 99564 22432
rect 99432 22392 99564 22420
rect 99432 22380 99438 22392
rect 99558 22380 99564 22392
rect 99616 22380 99622 22432
rect 1104 22330 1932 22352
rect 1104 22278 1322 22330
rect 1374 22278 1386 22330
rect 1438 22278 1932 22330
rect 1104 22256 1932 22278
rect 97980 22330 100832 22352
rect 97980 22278 98930 22330
rect 98982 22278 98994 22330
rect 99046 22278 99058 22330
rect 99110 22278 99122 22330
rect 99174 22278 99186 22330
rect 99238 22278 100832 22330
rect 97980 22256 100832 22278
rect 98457 22219 98515 22225
rect 98457 22185 98469 22219
rect 98503 22216 98515 22219
rect 99466 22216 99472 22228
rect 98503 22188 99472 22216
rect 98503 22185 98515 22188
rect 98457 22179 98515 22185
rect 99466 22176 99472 22188
rect 99524 22176 99530 22228
rect 97534 21904 97540 21956
rect 97592 21944 97598 21956
rect 98270 21944 98276 21956
rect 97592 21916 98276 21944
rect 97592 21904 97598 21916
rect 98270 21904 98276 21916
rect 98328 21904 98334 21956
rect 98489 21947 98547 21953
rect 98489 21913 98501 21947
rect 98535 21944 98547 21947
rect 98730 21944 98736 21956
rect 98535 21916 98736 21944
rect 98535 21913 98547 21916
rect 98489 21907 98547 21913
rect 98730 21904 98736 21916
rect 98788 21904 98794 21956
rect 98638 21836 98644 21888
rect 98696 21876 98702 21888
rect 99282 21876 99288 21888
rect 98696 21848 99288 21876
rect 98696 21836 98702 21848
rect 99282 21836 99288 21848
rect 99340 21836 99346 21888
rect 1104 21786 1932 21808
rect 1104 21734 1690 21786
rect 1742 21734 1754 21786
rect 1806 21734 1932 21786
rect 1104 21712 1932 21734
rect 97980 21786 100832 21808
rect 97980 21734 99666 21786
rect 99718 21734 99730 21786
rect 99782 21734 99794 21786
rect 99846 21734 99858 21786
rect 99910 21734 99922 21786
rect 99974 21734 100832 21786
rect 97980 21712 100832 21734
rect 1104 21242 1932 21264
rect 1104 21190 1322 21242
rect 1374 21190 1386 21242
rect 1438 21190 1932 21242
rect 1104 21168 1932 21190
rect 97980 21242 100832 21264
rect 97980 21190 98930 21242
rect 98982 21190 98994 21242
rect 99046 21190 99058 21242
rect 99110 21190 99122 21242
rect 99174 21190 99186 21242
rect 99238 21190 100832 21242
rect 97980 21168 100832 21190
rect 1104 20698 1932 20720
rect 1104 20646 1690 20698
rect 1742 20646 1754 20698
rect 1806 20646 1932 20698
rect 1104 20624 1932 20646
rect 97980 20698 100832 20720
rect 97980 20646 99666 20698
rect 99718 20646 99730 20698
rect 99782 20646 99794 20698
rect 99846 20646 99858 20698
rect 99910 20646 99922 20698
rect 99974 20646 100832 20698
rect 97980 20624 100832 20646
rect 1104 20154 1932 20176
rect 1104 20102 1322 20154
rect 1374 20102 1386 20154
rect 1438 20102 1932 20154
rect 1104 20080 1932 20102
rect 97980 20154 100832 20176
rect 97980 20102 98930 20154
rect 98982 20102 98994 20154
rect 99046 20102 99058 20154
rect 99110 20102 99122 20154
rect 99174 20102 99186 20154
rect 99238 20102 100832 20154
rect 97980 20080 100832 20102
rect 98822 19864 98828 19916
rect 98880 19904 98886 19916
rect 99837 19907 99895 19913
rect 99837 19904 99849 19907
rect 98880 19876 99849 19904
rect 98880 19864 98886 19876
rect 99837 19873 99849 19876
rect 99883 19873 99895 19907
rect 99837 19867 99895 19873
rect 100113 19907 100171 19913
rect 100113 19873 100125 19907
rect 100159 19904 100171 19907
rect 100202 19904 100208 19916
rect 100159 19876 100208 19904
rect 100159 19873 100171 19876
rect 100113 19867 100171 19873
rect 100202 19864 100208 19876
rect 100260 19864 100266 19916
rect 98454 19728 98460 19780
rect 98512 19768 98518 19780
rect 98512 19740 98670 19768
rect 98512 19728 98518 19740
rect 98362 19660 98368 19712
rect 98420 19660 98426 19712
rect 1104 19610 1932 19632
rect 1104 19558 1690 19610
rect 1742 19558 1754 19610
rect 1806 19558 1932 19610
rect 1104 19536 1932 19558
rect 97980 19610 100832 19632
rect 97980 19558 99666 19610
rect 99718 19558 99730 19610
rect 99782 19558 99794 19610
rect 99846 19558 99858 19610
rect 99910 19558 99922 19610
rect 99974 19558 100832 19610
rect 97980 19536 100832 19558
rect 98362 19252 98368 19304
rect 98420 19292 98426 19304
rect 99009 19295 99067 19301
rect 99009 19292 99021 19295
rect 98420 19264 99021 19292
rect 98420 19252 98426 19264
rect 99009 19261 99021 19264
rect 99055 19261 99067 19295
rect 99009 19255 99067 19261
rect 98454 19116 98460 19168
rect 98512 19116 98518 19168
rect 1104 19066 1932 19088
rect 1104 19014 1322 19066
rect 1374 19014 1386 19066
rect 1438 19014 1932 19066
rect 1104 18992 1932 19014
rect 97980 19066 100832 19088
rect 97980 19014 98930 19066
rect 98982 19014 98994 19066
rect 99046 19014 99058 19066
rect 99110 19014 99122 19066
rect 99174 19014 99186 19066
rect 99238 19014 100832 19066
rect 97980 18992 100832 19014
rect 1104 18522 1932 18544
rect 1104 18470 1690 18522
rect 1742 18470 1754 18522
rect 1806 18470 1932 18522
rect 1104 18448 1932 18470
rect 97980 18522 100832 18544
rect 97980 18470 99666 18522
rect 99718 18470 99730 18522
rect 99782 18470 99794 18522
rect 99846 18470 99858 18522
rect 99910 18470 99922 18522
rect 99974 18470 100832 18522
rect 97980 18448 100832 18470
rect 98454 18232 98460 18284
rect 98512 18232 98518 18284
rect 98549 18207 98607 18213
rect 98549 18173 98561 18207
rect 98595 18204 98607 18207
rect 98638 18204 98644 18216
rect 98595 18176 98644 18204
rect 98595 18173 98607 18176
rect 98549 18167 98607 18173
rect 98638 18164 98644 18176
rect 98696 18164 98702 18216
rect 98822 18164 98828 18216
rect 98880 18164 98886 18216
rect 1104 17978 1932 18000
rect 1104 17926 1322 17978
rect 1374 17926 1386 17978
rect 1438 17926 1932 17978
rect 1104 17904 1932 17926
rect 97980 17978 100832 18000
rect 97980 17926 98930 17978
rect 98982 17926 98994 17978
rect 99046 17926 99058 17978
rect 99110 17926 99122 17978
rect 99174 17926 99186 17978
rect 99238 17926 100832 17978
rect 97980 17904 100832 17926
rect 1104 17434 1932 17456
rect 1104 17382 1690 17434
rect 1742 17382 1754 17434
rect 1806 17382 1932 17434
rect 1104 17360 1932 17382
rect 97980 17434 100832 17456
rect 97980 17382 99666 17434
rect 99718 17382 99730 17434
rect 99782 17382 99794 17434
rect 99846 17382 99858 17434
rect 99910 17382 99922 17434
rect 99974 17382 100832 17434
rect 97980 17360 100832 17382
rect 1104 16890 1932 16912
rect 1104 16838 1322 16890
rect 1374 16838 1386 16890
rect 1438 16838 1932 16890
rect 1104 16816 1932 16838
rect 97980 16890 100832 16912
rect 97980 16838 98930 16890
rect 98982 16838 98994 16890
rect 99046 16838 99058 16890
rect 99110 16838 99122 16890
rect 99174 16838 99186 16890
rect 99238 16838 100832 16890
rect 97980 16816 100832 16838
rect 1104 16346 1932 16368
rect 1104 16294 1690 16346
rect 1742 16294 1754 16346
rect 1806 16294 1932 16346
rect 1104 16272 1932 16294
rect 97980 16346 100832 16368
rect 97980 16294 99666 16346
rect 99718 16294 99730 16346
rect 99782 16294 99794 16346
rect 99846 16294 99858 16346
rect 99910 16294 99922 16346
rect 99974 16294 100832 16346
rect 97980 16272 100832 16294
rect 1104 15802 1932 15824
rect 1104 15750 1322 15802
rect 1374 15750 1386 15802
rect 1438 15750 1932 15802
rect 1104 15728 1932 15750
rect 97980 15802 100832 15824
rect 97980 15750 98930 15802
rect 98982 15750 98994 15802
rect 99046 15750 99058 15802
rect 99110 15750 99122 15802
rect 99174 15750 99186 15802
rect 99238 15750 100832 15802
rect 97980 15728 100832 15750
rect 1104 15258 1932 15280
rect 1104 15206 1690 15258
rect 1742 15206 1754 15258
rect 1806 15206 1932 15258
rect 1104 15184 1932 15206
rect 97980 15258 100832 15280
rect 97980 15206 99666 15258
rect 99718 15206 99730 15258
rect 99782 15206 99794 15258
rect 99846 15206 99858 15258
rect 99910 15206 99922 15258
rect 99974 15206 100832 15258
rect 97980 15184 100832 15206
rect 1104 14714 1932 14736
rect 1104 14662 1322 14714
rect 1374 14662 1386 14714
rect 1438 14662 1932 14714
rect 1104 14640 1932 14662
rect 97980 14714 100832 14736
rect 97980 14662 98930 14714
rect 98982 14662 98994 14714
rect 99046 14662 99058 14714
rect 99110 14662 99122 14714
rect 99174 14662 99186 14714
rect 99238 14662 100832 14714
rect 97980 14640 100832 14662
rect 1104 14170 1932 14192
rect 1104 14118 1690 14170
rect 1742 14118 1754 14170
rect 1806 14118 1932 14170
rect 1104 14096 1932 14118
rect 97980 14170 100832 14192
rect 97980 14118 99666 14170
rect 99718 14118 99730 14170
rect 99782 14118 99794 14170
rect 99846 14118 99858 14170
rect 99910 14118 99922 14170
rect 99974 14118 100832 14170
rect 97980 14096 100832 14118
rect 1104 13626 1932 13648
rect 1104 13574 1322 13626
rect 1374 13574 1386 13626
rect 1438 13574 1932 13626
rect 1104 13552 1932 13574
rect 97980 13626 100832 13648
rect 97980 13574 98930 13626
rect 98982 13574 98994 13626
rect 99046 13574 99058 13626
rect 99110 13574 99122 13626
rect 99174 13574 99186 13626
rect 99238 13574 100832 13626
rect 97980 13552 100832 13574
rect 1104 13082 1932 13104
rect 1104 13030 1690 13082
rect 1742 13030 1754 13082
rect 1806 13030 1932 13082
rect 1104 13008 1932 13030
rect 97980 13082 100832 13104
rect 97980 13030 99666 13082
rect 99718 13030 99730 13082
rect 99782 13030 99794 13082
rect 99846 13030 99858 13082
rect 99910 13030 99922 13082
rect 99974 13030 100832 13082
rect 97980 13008 100832 13030
rect 1104 12538 1932 12560
rect 1104 12486 1322 12538
rect 1374 12486 1386 12538
rect 1438 12486 1932 12538
rect 1104 12464 1932 12486
rect 97980 12538 100832 12560
rect 97980 12486 98930 12538
rect 98982 12486 98994 12538
rect 99046 12486 99058 12538
rect 99110 12486 99122 12538
rect 99174 12486 99186 12538
rect 99238 12486 100832 12538
rect 97980 12464 100832 12486
rect 1104 11994 1932 12016
rect 1104 11942 1690 11994
rect 1742 11942 1754 11994
rect 1806 11942 1932 11994
rect 1104 11920 1932 11942
rect 97980 11994 100832 12016
rect 97980 11942 99666 11994
rect 99718 11942 99730 11994
rect 99782 11942 99794 11994
rect 99846 11942 99858 11994
rect 99910 11942 99922 11994
rect 99974 11942 100832 11994
rect 97980 11920 100832 11942
rect 1104 11450 1932 11472
rect 1104 11398 1322 11450
rect 1374 11398 1386 11450
rect 1438 11398 1932 11450
rect 1104 11376 1932 11398
rect 97980 11450 100832 11472
rect 97980 11398 98930 11450
rect 98982 11398 98994 11450
rect 99046 11398 99058 11450
rect 99110 11398 99122 11450
rect 99174 11398 99186 11450
rect 99238 11398 100832 11450
rect 97980 11376 100832 11398
rect 1104 10906 1932 10928
rect 1104 10854 1690 10906
rect 1742 10854 1754 10906
rect 1806 10854 1932 10906
rect 1104 10832 1932 10854
rect 97980 10906 100832 10928
rect 97980 10854 99666 10906
rect 99718 10854 99730 10906
rect 99782 10854 99794 10906
rect 99846 10854 99858 10906
rect 99910 10854 99922 10906
rect 99974 10854 100832 10906
rect 97980 10832 100832 10854
rect 1104 10362 1932 10384
rect 1104 10310 1322 10362
rect 1374 10310 1386 10362
rect 1438 10310 1932 10362
rect 1104 10288 1932 10310
rect 97980 10362 100832 10384
rect 97980 10310 98930 10362
rect 98982 10310 98994 10362
rect 99046 10310 99058 10362
rect 99110 10310 99122 10362
rect 99174 10310 99186 10362
rect 99238 10310 100832 10362
rect 97980 10288 100832 10310
rect 1104 9818 1932 9840
rect 1104 9766 1690 9818
rect 1742 9766 1754 9818
rect 1806 9766 1932 9818
rect 1104 9744 1932 9766
rect 97980 9818 100832 9840
rect 97980 9766 99666 9818
rect 99718 9766 99730 9818
rect 99782 9766 99794 9818
rect 99846 9766 99858 9818
rect 99910 9766 99922 9818
rect 99974 9766 100832 9818
rect 97980 9744 100832 9766
rect 1104 9274 1932 9296
rect 1104 9222 1322 9274
rect 1374 9222 1386 9274
rect 1438 9222 1932 9274
rect 1104 9200 1932 9222
rect 97980 9274 100832 9296
rect 97980 9222 98930 9274
rect 98982 9222 98994 9274
rect 99046 9222 99058 9274
rect 99110 9222 99122 9274
rect 99174 9222 99186 9274
rect 99238 9222 100832 9274
rect 97980 9200 100832 9222
rect 1104 8730 1932 8752
rect 1104 8678 1690 8730
rect 1742 8678 1754 8730
rect 1806 8678 1932 8730
rect 1104 8656 1932 8678
rect 97980 8730 100832 8752
rect 97980 8678 99666 8730
rect 99718 8678 99730 8730
rect 99782 8678 99794 8730
rect 99846 8678 99858 8730
rect 99910 8678 99922 8730
rect 99974 8678 100832 8730
rect 97980 8656 100832 8678
rect 1104 8186 1932 8208
rect 1104 8134 1322 8186
rect 1374 8134 1386 8186
rect 1438 8134 1932 8186
rect 1104 8112 1932 8134
rect 97980 8186 100832 8208
rect 97980 8134 98930 8186
rect 98982 8134 98994 8186
rect 99046 8134 99058 8186
rect 99110 8134 99122 8186
rect 99174 8134 99186 8186
rect 99238 8134 100832 8186
rect 97980 8112 100832 8134
rect 1104 7642 1932 7664
rect 1104 7590 1690 7642
rect 1742 7590 1754 7642
rect 1806 7590 1932 7642
rect 1104 7568 1932 7590
rect 97980 7642 100832 7664
rect 97980 7590 99666 7642
rect 99718 7590 99730 7642
rect 99782 7590 99794 7642
rect 99846 7590 99858 7642
rect 99910 7590 99922 7642
rect 99974 7590 100832 7642
rect 97980 7568 100832 7590
rect 1104 7098 1932 7120
rect 1104 7046 1322 7098
rect 1374 7046 1386 7098
rect 1438 7046 1932 7098
rect 1104 7024 1932 7046
rect 97980 7098 100832 7120
rect 97980 7046 98930 7098
rect 98982 7046 98994 7098
rect 99046 7046 99058 7098
rect 99110 7046 99122 7098
rect 99174 7046 99186 7098
rect 99238 7046 100832 7098
rect 97980 7024 100832 7046
rect 1104 6554 1932 6576
rect 1104 6502 1690 6554
rect 1742 6502 1754 6554
rect 1806 6502 1932 6554
rect 1104 6480 1932 6502
rect 97980 6554 100832 6576
rect 97980 6502 99666 6554
rect 99718 6502 99730 6554
rect 99782 6502 99794 6554
rect 99846 6502 99858 6554
rect 99910 6502 99922 6554
rect 99974 6502 100832 6554
rect 97980 6480 100832 6502
rect 1104 6010 1932 6032
rect 1104 5958 1322 6010
rect 1374 5958 1386 6010
rect 1438 5958 1932 6010
rect 1104 5936 1932 5958
rect 97980 6010 100832 6032
rect 97980 5958 98930 6010
rect 98982 5958 98994 6010
rect 99046 5958 99058 6010
rect 99110 5958 99122 6010
rect 99174 5958 99186 6010
rect 99238 5958 100832 6010
rect 97980 5936 100832 5958
rect 1104 5466 1932 5488
rect 1104 5414 1690 5466
rect 1742 5414 1754 5466
rect 1806 5414 1932 5466
rect 1104 5392 1932 5414
rect 97980 5466 100832 5488
rect 97980 5414 99666 5466
rect 99718 5414 99730 5466
rect 99782 5414 99794 5466
rect 99846 5414 99858 5466
rect 99910 5414 99922 5466
rect 99974 5414 100832 5466
rect 97980 5392 100832 5414
rect 1104 4922 1932 4944
rect 1104 4870 1322 4922
rect 1374 4870 1386 4922
rect 1438 4870 1932 4922
rect 1104 4848 1932 4870
rect 97980 4922 100832 4944
rect 97980 4870 98930 4922
rect 98982 4870 98994 4922
rect 99046 4870 99058 4922
rect 99110 4870 99122 4922
rect 99174 4870 99186 4922
rect 99238 4870 100832 4922
rect 97980 4848 100832 4870
rect 1104 4378 1932 4400
rect 1104 4326 1690 4378
rect 1742 4326 1754 4378
rect 1806 4326 1932 4378
rect 1104 4304 1932 4326
rect 97980 4378 100832 4400
rect 97980 4326 99666 4378
rect 99718 4326 99730 4378
rect 99782 4326 99794 4378
rect 99846 4326 99858 4378
rect 99910 4326 99922 4378
rect 99974 4326 100832 4378
rect 97980 4304 100832 4326
rect 1104 3834 1932 3856
rect 1104 3782 1322 3834
rect 1374 3782 1386 3834
rect 1438 3782 1932 3834
rect 1104 3760 1932 3782
rect 97980 3834 100832 3856
rect 97980 3782 98930 3834
rect 98982 3782 98994 3834
rect 99046 3782 99058 3834
rect 99110 3782 99122 3834
rect 99174 3782 99186 3834
rect 99238 3782 100832 3834
rect 97980 3760 100832 3782
rect 1104 3290 1932 3312
rect 1104 3238 1690 3290
rect 1742 3238 1754 3290
rect 1806 3238 1932 3290
rect 1104 3216 1932 3238
rect 97980 3290 100832 3312
rect 97980 3238 99666 3290
rect 99718 3238 99730 3290
rect 99782 3238 99794 3290
rect 99846 3238 99858 3290
rect 99910 3238 99922 3290
rect 99974 3238 100832 3290
rect 97980 3216 100832 3238
rect 1104 2746 1932 2768
rect 1104 2694 1322 2746
rect 1374 2694 1386 2746
rect 1438 2694 1932 2746
rect 1104 2672 1932 2694
rect 97980 2746 100832 2768
rect 97980 2694 98930 2746
rect 98982 2694 98994 2746
rect 99046 2694 99058 2746
rect 99110 2694 99122 2746
rect 99174 2694 99186 2746
rect 99238 2694 100832 2746
rect 97980 2672 100832 2694
rect 1104 2202 1932 2224
rect 1104 2150 1690 2202
rect 1742 2150 1754 2202
rect 1806 2150 1932 2202
rect 1104 2128 1932 2150
rect 97980 2202 100832 2224
rect 97980 2150 99666 2202
rect 99718 2150 99730 2202
rect 99782 2150 99794 2202
rect 99846 2150 99858 2202
rect 99910 2150 99922 2202
rect 99974 2150 100832 2202
rect 97980 2128 100832 2150
<< via1 >>
rect 4214 101702 4266 101754
rect 4278 101702 4330 101754
rect 4342 101702 4394 101754
rect 4406 101702 4458 101754
rect 4470 101702 4522 101754
rect 34934 101702 34986 101754
rect 34998 101702 35050 101754
rect 35062 101702 35114 101754
rect 35126 101702 35178 101754
rect 35190 101702 35242 101754
rect 65654 101702 65706 101754
rect 65718 101702 65770 101754
rect 65782 101702 65834 101754
rect 65846 101702 65898 101754
rect 65910 101702 65962 101754
rect 96374 101702 96426 101754
rect 96438 101702 96490 101754
rect 96502 101702 96554 101754
rect 96566 101702 96618 101754
rect 96630 101702 96682 101754
rect 43352 101643 43404 101652
rect 43352 101609 43361 101643
rect 43361 101609 43395 101643
rect 43395 101609 43404 101643
rect 43352 101600 43404 101609
rect 45284 101643 45336 101652
rect 45284 101609 45293 101643
rect 45293 101609 45327 101643
rect 45327 101609 45336 101643
rect 45284 101600 45336 101609
rect 47952 101643 48004 101652
rect 47952 101609 47961 101643
rect 47961 101609 47995 101643
rect 47995 101609 48004 101643
rect 47952 101600 48004 101609
rect 49516 101600 49568 101652
rect 50988 101600 51040 101652
rect 53012 101643 53064 101652
rect 53012 101609 53021 101643
rect 53021 101609 53055 101643
rect 53055 101609 53064 101643
rect 53012 101600 53064 101609
rect 55680 101643 55732 101652
rect 55680 101609 55689 101643
rect 55689 101609 55723 101643
rect 55723 101609 55732 101643
rect 55680 101600 55732 101609
rect 57612 101643 57664 101652
rect 57612 101609 57621 101643
rect 57621 101609 57655 101643
rect 57655 101609 57664 101643
rect 57612 101600 57664 101609
rect 58808 101643 58860 101652
rect 58808 101609 58817 101643
rect 58817 101609 58851 101643
rect 58851 101609 58860 101643
rect 58808 101600 58860 101609
rect 43536 101439 43588 101448
rect 43536 101405 43545 101439
rect 43545 101405 43579 101439
rect 43579 101405 43588 101439
rect 43536 101396 43588 101405
rect 45376 101396 45428 101448
rect 47492 101396 47544 101448
rect 49700 101439 49752 101448
rect 49700 101405 49709 101439
rect 49709 101405 49743 101439
rect 49743 101405 49752 101439
rect 49700 101396 49752 101405
rect 51172 101396 51224 101448
rect 53104 101396 53156 101448
rect 55128 101396 55180 101448
rect 57336 101396 57388 101448
rect 59176 101396 59228 101448
rect 4874 101158 4926 101210
rect 4938 101158 4990 101210
rect 5002 101158 5054 101210
rect 5066 101158 5118 101210
rect 5130 101158 5182 101210
rect 35594 101158 35646 101210
rect 35658 101158 35710 101210
rect 35722 101158 35774 101210
rect 35786 101158 35838 101210
rect 35850 101158 35902 101210
rect 66314 101158 66366 101210
rect 66378 101158 66430 101210
rect 66442 101158 66494 101210
rect 66506 101158 66558 101210
rect 66570 101158 66622 101210
rect 97034 101158 97086 101210
rect 97098 101158 97150 101210
rect 97162 101158 97214 101210
rect 97226 101158 97278 101210
rect 97290 101158 97342 101210
rect 4214 100614 4266 100666
rect 4278 100614 4330 100666
rect 4342 100614 4394 100666
rect 4406 100614 4458 100666
rect 4470 100614 4522 100666
rect 34934 100614 34986 100666
rect 34998 100614 35050 100666
rect 35062 100614 35114 100666
rect 35126 100614 35178 100666
rect 35190 100614 35242 100666
rect 65654 100614 65706 100666
rect 65718 100614 65770 100666
rect 65782 100614 65834 100666
rect 65846 100614 65898 100666
rect 65910 100614 65962 100666
rect 96374 100614 96426 100666
rect 96438 100614 96490 100666
rect 96502 100614 96554 100666
rect 96566 100614 96618 100666
rect 96630 100614 96682 100666
rect 4874 100070 4926 100122
rect 4938 100070 4990 100122
rect 5002 100070 5054 100122
rect 5066 100070 5118 100122
rect 5130 100070 5182 100122
rect 35594 100070 35646 100122
rect 35658 100070 35710 100122
rect 35722 100070 35774 100122
rect 35786 100070 35838 100122
rect 35850 100070 35902 100122
rect 66314 100070 66366 100122
rect 66378 100070 66430 100122
rect 66442 100070 66494 100122
rect 66506 100070 66558 100122
rect 66570 100070 66622 100122
rect 97034 100070 97086 100122
rect 97098 100070 97150 100122
rect 97162 100070 97214 100122
rect 97226 100070 97278 100122
rect 97290 100070 97342 100122
rect 4214 99526 4266 99578
rect 4278 99526 4330 99578
rect 4342 99526 4394 99578
rect 4406 99526 4458 99578
rect 4470 99526 4522 99578
rect 34934 99526 34986 99578
rect 34998 99526 35050 99578
rect 35062 99526 35114 99578
rect 35126 99526 35178 99578
rect 35190 99526 35242 99578
rect 65654 99526 65706 99578
rect 65718 99526 65770 99578
rect 65782 99526 65834 99578
rect 65846 99526 65898 99578
rect 65910 99526 65962 99578
rect 96374 99526 96426 99578
rect 96438 99526 96490 99578
rect 96502 99526 96554 99578
rect 96566 99526 96618 99578
rect 96630 99526 96682 99578
rect 4874 98982 4926 99034
rect 4938 98982 4990 99034
rect 5002 98982 5054 99034
rect 5066 98982 5118 99034
rect 5130 98982 5182 99034
rect 35594 98982 35646 99034
rect 35658 98982 35710 99034
rect 35722 98982 35774 99034
rect 35786 98982 35838 99034
rect 35850 98982 35902 99034
rect 66314 98982 66366 99034
rect 66378 98982 66430 99034
rect 66442 98982 66494 99034
rect 66506 98982 66558 99034
rect 66570 98982 66622 99034
rect 97034 98982 97086 99034
rect 97098 98982 97150 99034
rect 97162 98982 97214 99034
rect 97226 98982 97278 99034
rect 97290 98982 97342 99034
rect 4214 98438 4266 98490
rect 4278 98438 4330 98490
rect 4342 98438 4394 98490
rect 4406 98438 4458 98490
rect 4470 98438 4522 98490
rect 34934 98438 34986 98490
rect 34998 98438 35050 98490
rect 35062 98438 35114 98490
rect 35126 98438 35178 98490
rect 35190 98438 35242 98490
rect 65654 98438 65706 98490
rect 65718 98438 65770 98490
rect 65782 98438 65834 98490
rect 65846 98438 65898 98490
rect 65910 98438 65962 98490
rect 96374 98438 96426 98490
rect 96438 98438 96490 98490
rect 96502 98438 96554 98490
rect 96566 98438 96618 98490
rect 96630 98438 96682 98490
rect 4874 97894 4926 97946
rect 4938 97894 4990 97946
rect 5002 97894 5054 97946
rect 5066 97894 5118 97946
rect 5130 97894 5182 97946
rect 35594 97894 35646 97946
rect 35658 97894 35710 97946
rect 35722 97894 35774 97946
rect 35786 97894 35838 97946
rect 35850 97894 35902 97946
rect 66314 97894 66366 97946
rect 66378 97894 66430 97946
rect 66442 97894 66494 97946
rect 66506 97894 66558 97946
rect 66570 97894 66622 97946
rect 97034 97894 97086 97946
rect 97098 97894 97150 97946
rect 97162 97894 97214 97946
rect 97226 97894 97278 97946
rect 97290 97894 97342 97946
rect 4214 97350 4266 97402
rect 4278 97350 4330 97402
rect 4342 97350 4394 97402
rect 4406 97350 4458 97402
rect 4470 97350 4522 97402
rect 34934 97350 34986 97402
rect 34998 97350 35050 97402
rect 35062 97350 35114 97402
rect 35126 97350 35178 97402
rect 35190 97350 35242 97402
rect 65654 97350 65706 97402
rect 65718 97350 65770 97402
rect 65782 97350 65834 97402
rect 65846 97350 65898 97402
rect 65910 97350 65962 97402
rect 96374 97350 96426 97402
rect 96438 97350 96490 97402
rect 96502 97350 96554 97402
rect 96566 97350 96618 97402
rect 96630 97350 96682 97402
rect 4874 96806 4926 96858
rect 4938 96806 4990 96858
rect 5002 96806 5054 96858
rect 5066 96806 5118 96858
rect 5130 96806 5182 96858
rect 35594 96806 35646 96858
rect 35658 96806 35710 96858
rect 35722 96806 35774 96858
rect 35786 96806 35838 96858
rect 35850 96806 35902 96858
rect 66314 96806 66366 96858
rect 66378 96806 66430 96858
rect 66442 96806 66494 96858
rect 66506 96806 66558 96858
rect 66570 96806 66622 96858
rect 97034 96806 97086 96858
rect 97098 96806 97150 96858
rect 97162 96806 97214 96858
rect 97226 96806 97278 96858
rect 97290 96806 97342 96858
rect 4214 96262 4266 96314
rect 4278 96262 4330 96314
rect 4342 96262 4394 96314
rect 4406 96262 4458 96314
rect 4470 96262 4522 96314
rect 34934 96262 34986 96314
rect 34998 96262 35050 96314
rect 35062 96262 35114 96314
rect 35126 96262 35178 96314
rect 35190 96262 35242 96314
rect 65654 96262 65706 96314
rect 65718 96262 65770 96314
rect 65782 96262 65834 96314
rect 65846 96262 65898 96314
rect 65910 96262 65962 96314
rect 96374 96262 96426 96314
rect 96438 96262 96490 96314
rect 96502 96262 96554 96314
rect 96566 96262 96618 96314
rect 96630 96262 96682 96314
rect 4874 95718 4926 95770
rect 4938 95718 4990 95770
rect 5002 95718 5054 95770
rect 5066 95718 5118 95770
rect 5130 95718 5182 95770
rect 35594 95718 35646 95770
rect 35658 95718 35710 95770
rect 35722 95718 35774 95770
rect 35786 95718 35838 95770
rect 35850 95718 35902 95770
rect 66314 95718 66366 95770
rect 66378 95718 66430 95770
rect 66442 95718 66494 95770
rect 66506 95718 66558 95770
rect 66570 95718 66622 95770
rect 97034 95718 97086 95770
rect 97098 95718 97150 95770
rect 97162 95718 97214 95770
rect 97226 95718 97278 95770
rect 97290 95718 97342 95770
rect 4214 95174 4266 95226
rect 4278 95174 4330 95226
rect 4342 95174 4394 95226
rect 4406 95174 4458 95226
rect 4470 95174 4522 95226
rect 34934 95174 34986 95226
rect 34998 95174 35050 95226
rect 35062 95174 35114 95226
rect 35126 95174 35178 95226
rect 35190 95174 35242 95226
rect 65654 95174 65706 95226
rect 65718 95174 65770 95226
rect 65782 95174 65834 95226
rect 65846 95174 65898 95226
rect 65910 95174 65962 95226
rect 96374 95174 96426 95226
rect 96438 95174 96490 95226
rect 96502 95174 96554 95226
rect 96566 95174 96618 95226
rect 96630 95174 96682 95226
rect 4874 94630 4926 94682
rect 4938 94630 4990 94682
rect 5002 94630 5054 94682
rect 5066 94630 5118 94682
rect 5130 94630 5182 94682
rect 35594 94630 35646 94682
rect 35658 94630 35710 94682
rect 35722 94630 35774 94682
rect 35786 94630 35838 94682
rect 35850 94630 35902 94682
rect 66314 94630 66366 94682
rect 66378 94630 66430 94682
rect 66442 94630 66494 94682
rect 66506 94630 66558 94682
rect 66570 94630 66622 94682
rect 97034 94630 97086 94682
rect 97098 94630 97150 94682
rect 97162 94630 97214 94682
rect 97226 94630 97278 94682
rect 97290 94630 97342 94682
rect 4214 94086 4266 94138
rect 4278 94086 4330 94138
rect 4342 94086 4394 94138
rect 4406 94086 4458 94138
rect 4470 94086 4522 94138
rect 34934 94086 34986 94138
rect 34998 94086 35050 94138
rect 35062 94086 35114 94138
rect 35126 94086 35178 94138
rect 35190 94086 35242 94138
rect 65654 94086 65706 94138
rect 65718 94086 65770 94138
rect 65782 94086 65834 94138
rect 65846 94086 65898 94138
rect 65910 94086 65962 94138
rect 96374 94086 96426 94138
rect 96438 94086 96490 94138
rect 96502 94086 96554 94138
rect 96566 94086 96618 94138
rect 96630 94086 96682 94138
rect 4874 93542 4926 93594
rect 4938 93542 4990 93594
rect 5002 93542 5054 93594
rect 5066 93542 5118 93594
rect 5130 93542 5182 93594
rect 35594 93542 35646 93594
rect 35658 93542 35710 93594
rect 35722 93542 35774 93594
rect 35786 93542 35838 93594
rect 35850 93542 35902 93594
rect 66314 93542 66366 93594
rect 66378 93542 66430 93594
rect 66442 93542 66494 93594
rect 66506 93542 66558 93594
rect 66570 93542 66622 93594
rect 97034 93542 97086 93594
rect 97098 93542 97150 93594
rect 97162 93542 97214 93594
rect 97226 93542 97278 93594
rect 97290 93542 97342 93594
rect 4214 92998 4266 93050
rect 4278 92998 4330 93050
rect 4342 92998 4394 93050
rect 4406 92998 4458 93050
rect 4470 92998 4522 93050
rect 34934 92998 34986 93050
rect 34998 92998 35050 93050
rect 35062 92998 35114 93050
rect 35126 92998 35178 93050
rect 35190 92998 35242 93050
rect 65654 92998 65706 93050
rect 65718 92998 65770 93050
rect 65782 92998 65834 93050
rect 65846 92998 65898 93050
rect 65910 92998 65962 93050
rect 96374 92998 96426 93050
rect 96438 92998 96490 93050
rect 96502 92998 96554 93050
rect 96566 92998 96618 93050
rect 96630 92998 96682 93050
rect 4874 92454 4926 92506
rect 4938 92454 4990 92506
rect 5002 92454 5054 92506
rect 5066 92454 5118 92506
rect 5130 92454 5182 92506
rect 35594 92454 35646 92506
rect 35658 92454 35710 92506
rect 35722 92454 35774 92506
rect 35786 92454 35838 92506
rect 35850 92454 35902 92506
rect 66314 92454 66366 92506
rect 66378 92454 66430 92506
rect 66442 92454 66494 92506
rect 66506 92454 66558 92506
rect 66570 92454 66622 92506
rect 97034 92454 97086 92506
rect 97098 92454 97150 92506
rect 97162 92454 97214 92506
rect 97226 92454 97278 92506
rect 97290 92454 97342 92506
rect 4214 91910 4266 91962
rect 4278 91910 4330 91962
rect 4342 91910 4394 91962
rect 4406 91910 4458 91962
rect 4470 91910 4522 91962
rect 34934 91910 34986 91962
rect 34998 91910 35050 91962
rect 35062 91910 35114 91962
rect 35126 91910 35178 91962
rect 35190 91910 35242 91962
rect 65654 91910 65706 91962
rect 65718 91910 65770 91962
rect 65782 91910 65834 91962
rect 65846 91910 65898 91962
rect 65910 91910 65962 91962
rect 96374 91910 96426 91962
rect 96438 91910 96490 91962
rect 96502 91910 96554 91962
rect 96566 91910 96618 91962
rect 96630 91910 96682 91962
rect 4874 91366 4926 91418
rect 4938 91366 4990 91418
rect 5002 91366 5054 91418
rect 5066 91366 5118 91418
rect 5130 91366 5182 91418
rect 35594 91366 35646 91418
rect 35658 91366 35710 91418
rect 35722 91366 35774 91418
rect 35786 91366 35838 91418
rect 35850 91366 35902 91418
rect 66314 91366 66366 91418
rect 66378 91366 66430 91418
rect 66442 91366 66494 91418
rect 66506 91366 66558 91418
rect 66570 91366 66622 91418
rect 97034 91366 97086 91418
rect 97098 91366 97150 91418
rect 97162 91366 97214 91418
rect 97226 91366 97278 91418
rect 97290 91366 97342 91418
rect 4214 90822 4266 90874
rect 4278 90822 4330 90874
rect 4342 90822 4394 90874
rect 4406 90822 4458 90874
rect 4470 90822 4522 90874
rect 34934 90822 34986 90874
rect 34998 90822 35050 90874
rect 35062 90822 35114 90874
rect 35126 90822 35178 90874
rect 35190 90822 35242 90874
rect 65654 90822 65706 90874
rect 65718 90822 65770 90874
rect 65782 90822 65834 90874
rect 65846 90822 65898 90874
rect 65910 90822 65962 90874
rect 96374 90822 96426 90874
rect 96438 90822 96490 90874
rect 96502 90822 96554 90874
rect 96566 90822 96618 90874
rect 96630 90822 96682 90874
rect 4874 90278 4926 90330
rect 4938 90278 4990 90330
rect 5002 90278 5054 90330
rect 5066 90278 5118 90330
rect 5130 90278 5182 90330
rect 35594 90278 35646 90330
rect 35658 90278 35710 90330
rect 35722 90278 35774 90330
rect 35786 90278 35838 90330
rect 35850 90278 35902 90330
rect 66314 90278 66366 90330
rect 66378 90278 66430 90330
rect 66442 90278 66494 90330
rect 66506 90278 66558 90330
rect 66570 90278 66622 90330
rect 97034 90278 97086 90330
rect 97098 90278 97150 90330
rect 97162 90278 97214 90330
rect 97226 90278 97278 90330
rect 97290 90278 97342 90330
rect 4214 89734 4266 89786
rect 4278 89734 4330 89786
rect 4342 89734 4394 89786
rect 4406 89734 4458 89786
rect 4470 89734 4522 89786
rect 34934 89734 34986 89786
rect 34998 89734 35050 89786
rect 35062 89734 35114 89786
rect 35126 89734 35178 89786
rect 35190 89734 35242 89786
rect 65654 89734 65706 89786
rect 65718 89734 65770 89786
rect 65782 89734 65834 89786
rect 65846 89734 65898 89786
rect 65910 89734 65962 89786
rect 96374 89734 96426 89786
rect 96438 89734 96490 89786
rect 96502 89734 96554 89786
rect 96566 89734 96618 89786
rect 96630 89734 96682 89786
rect 4874 89190 4926 89242
rect 4938 89190 4990 89242
rect 5002 89190 5054 89242
rect 5066 89190 5118 89242
rect 5130 89190 5182 89242
rect 35594 89190 35646 89242
rect 35658 89190 35710 89242
rect 35722 89190 35774 89242
rect 35786 89190 35838 89242
rect 35850 89190 35902 89242
rect 66314 89190 66366 89242
rect 66378 89190 66430 89242
rect 66442 89190 66494 89242
rect 66506 89190 66558 89242
rect 66570 89190 66622 89242
rect 97034 89190 97086 89242
rect 97098 89190 97150 89242
rect 97162 89190 97214 89242
rect 97226 89190 97278 89242
rect 97290 89190 97342 89242
rect 4214 88646 4266 88698
rect 4278 88646 4330 88698
rect 4342 88646 4394 88698
rect 4406 88646 4458 88698
rect 4470 88646 4522 88698
rect 34934 88646 34986 88698
rect 34998 88646 35050 88698
rect 35062 88646 35114 88698
rect 35126 88646 35178 88698
rect 35190 88646 35242 88698
rect 65654 88646 65706 88698
rect 65718 88646 65770 88698
rect 65782 88646 65834 88698
rect 65846 88646 65898 88698
rect 65910 88646 65962 88698
rect 96374 88646 96426 88698
rect 96438 88646 96490 88698
rect 96502 88646 96554 88698
rect 96566 88646 96618 88698
rect 96630 88646 96682 88698
rect 4874 88102 4926 88154
rect 4938 88102 4990 88154
rect 5002 88102 5054 88154
rect 5066 88102 5118 88154
rect 5130 88102 5182 88154
rect 35594 88102 35646 88154
rect 35658 88102 35710 88154
rect 35722 88102 35774 88154
rect 35786 88102 35838 88154
rect 35850 88102 35902 88154
rect 66314 88102 66366 88154
rect 66378 88102 66430 88154
rect 66442 88102 66494 88154
rect 66506 88102 66558 88154
rect 66570 88102 66622 88154
rect 97034 88102 97086 88154
rect 97098 88102 97150 88154
rect 97162 88102 97214 88154
rect 97226 88102 97278 88154
rect 97290 88102 97342 88154
rect 4214 87558 4266 87610
rect 4278 87558 4330 87610
rect 4342 87558 4394 87610
rect 4406 87558 4458 87610
rect 4470 87558 4522 87610
rect 34934 87558 34986 87610
rect 34998 87558 35050 87610
rect 35062 87558 35114 87610
rect 35126 87558 35178 87610
rect 35190 87558 35242 87610
rect 65654 87558 65706 87610
rect 65718 87558 65770 87610
rect 65782 87558 65834 87610
rect 65846 87558 65898 87610
rect 65910 87558 65962 87610
rect 96374 87558 96426 87610
rect 96438 87558 96490 87610
rect 96502 87558 96554 87610
rect 96566 87558 96618 87610
rect 96630 87558 96682 87610
rect 4874 87014 4926 87066
rect 4938 87014 4990 87066
rect 5002 87014 5054 87066
rect 5066 87014 5118 87066
rect 5130 87014 5182 87066
rect 35594 87014 35646 87066
rect 35658 87014 35710 87066
rect 35722 87014 35774 87066
rect 35786 87014 35838 87066
rect 35850 87014 35902 87066
rect 66314 87014 66366 87066
rect 66378 87014 66430 87066
rect 66442 87014 66494 87066
rect 66506 87014 66558 87066
rect 66570 87014 66622 87066
rect 97034 87014 97086 87066
rect 97098 87014 97150 87066
rect 97162 87014 97214 87066
rect 97226 87014 97278 87066
rect 97290 87014 97342 87066
rect 4214 86470 4266 86522
rect 4278 86470 4330 86522
rect 4342 86470 4394 86522
rect 4406 86470 4458 86522
rect 4470 86470 4522 86522
rect 34934 86470 34986 86522
rect 34998 86470 35050 86522
rect 35062 86470 35114 86522
rect 35126 86470 35178 86522
rect 35190 86470 35242 86522
rect 65654 86470 65706 86522
rect 65718 86470 65770 86522
rect 65782 86470 65834 86522
rect 65846 86470 65898 86522
rect 65910 86470 65962 86522
rect 96374 86470 96426 86522
rect 96438 86470 96490 86522
rect 96502 86470 96554 86522
rect 96566 86470 96618 86522
rect 96630 86470 96682 86522
rect 4874 85926 4926 85978
rect 4938 85926 4990 85978
rect 5002 85926 5054 85978
rect 5066 85926 5118 85978
rect 5130 85926 5182 85978
rect 35594 85926 35646 85978
rect 35658 85926 35710 85978
rect 35722 85926 35774 85978
rect 35786 85926 35838 85978
rect 35850 85926 35902 85978
rect 66314 85926 66366 85978
rect 66378 85926 66430 85978
rect 66442 85926 66494 85978
rect 66506 85926 66558 85978
rect 66570 85926 66622 85978
rect 97034 85926 97086 85978
rect 97098 85926 97150 85978
rect 97162 85926 97214 85978
rect 97226 85926 97278 85978
rect 97290 85926 97342 85978
rect 4214 85382 4266 85434
rect 4278 85382 4330 85434
rect 4342 85382 4394 85434
rect 4406 85382 4458 85434
rect 4470 85382 4522 85434
rect 34934 85382 34986 85434
rect 34998 85382 35050 85434
rect 35062 85382 35114 85434
rect 35126 85382 35178 85434
rect 35190 85382 35242 85434
rect 65654 85382 65706 85434
rect 65718 85382 65770 85434
rect 65782 85382 65834 85434
rect 65846 85382 65898 85434
rect 65910 85382 65962 85434
rect 96374 85382 96426 85434
rect 96438 85382 96490 85434
rect 96502 85382 96554 85434
rect 96566 85382 96618 85434
rect 96630 85382 96682 85434
rect 4874 84838 4926 84890
rect 4938 84838 4990 84890
rect 5002 84838 5054 84890
rect 5066 84838 5118 84890
rect 5130 84838 5182 84890
rect 35594 84838 35646 84890
rect 35658 84838 35710 84890
rect 35722 84838 35774 84890
rect 35786 84838 35838 84890
rect 35850 84838 35902 84890
rect 66314 84838 66366 84890
rect 66378 84838 66430 84890
rect 66442 84838 66494 84890
rect 66506 84838 66558 84890
rect 66570 84838 66622 84890
rect 97034 84838 97086 84890
rect 97098 84838 97150 84890
rect 97162 84838 97214 84890
rect 97226 84838 97278 84890
rect 97290 84838 97342 84890
rect 4214 84294 4266 84346
rect 4278 84294 4330 84346
rect 4342 84294 4394 84346
rect 4406 84294 4458 84346
rect 4470 84294 4522 84346
rect 34934 84294 34986 84346
rect 34998 84294 35050 84346
rect 35062 84294 35114 84346
rect 35126 84294 35178 84346
rect 35190 84294 35242 84346
rect 65654 84294 65706 84346
rect 65718 84294 65770 84346
rect 65782 84294 65834 84346
rect 65846 84294 65898 84346
rect 65910 84294 65962 84346
rect 96374 84294 96426 84346
rect 96438 84294 96490 84346
rect 96502 84294 96554 84346
rect 96566 84294 96618 84346
rect 96630 84294 96682 84346
rect 4874 83750 4926 83802
rect 4938 83750 4990 83802
rect 5002 83750 5054 83802
rect 5066 83750 5118 83802
rect 5130 83750 5182 83802
rect 35594 83750 35646 83802
rect 35658 83750 35710 83802
rect 35722 83750 35774 83802
rect 35786 83750 35838 83802
rect 35850 83750 35902 83802
rect 66314 83750 66366 83802
rect 66378 83750 66430 83802
rect 66442 83750 66494 83802
rect 66506 83750 66558 83802
rect 66570 83750 66622 83802
rect 97034 83750 97086 83802
rect 97098 83750 97150 83802
rect 97162 83750 97214 83802
rect 97226 83750 97278 83802
rect 97290 83750 97342 83802
rect 4214 83206 4266 83258
rect 4278 83206 4330 83258
rect 4342 83206 4394 83258
rect 4406 83206 4458 83258
rect 4470 83206 4522 83258
rect 34934 83206 34986 83258
rect 34998 83206 35050 83258
rect 35062 83206 35114 83258
rect 35126 83206 35178 83258
rect 35190 83206 35242 83258
rect 65654 83206 65706 83258
rect 65718 83206 65770 83258
rect 65782 83206 65834 83258
rect 65846 83206 65898 83258
rect 65910 83206 65962 83258
rect 96374 83206 96426 83258
rect 96438 83206 96490 83258
rect 96502 83206 96554 83258
rect 96566 83206 96618 83258
rect 96630 83206 96682 83258
rect 4874 82662 4926 82714
rect 4938 82662 4990 82714
rect 5002 82662 5054 82714
rect 5066 82662 5118 82714
rect 5130 82662 5182 82714
rect 35594 82662 35646 82714
rect 35658 82662 35710 82714
rect 35722 82662 35774 82714
rect 35786 82662 35838 82714
rect 35850 82662 35902 82714
rect 66314 82662 66366 82714
rect 66378 82662 66430 82714
rect 66442 82662 66494 82714
rect 66506 82662 66558 82714
rect 66570 82662 66622 82714
rect 97034 82662 97086 82714
rect 97098 82662 97150 82714
rect 97162 82662 97214 82714
rect 97226 82662 97278 82714
rect 97290 82662 97342 82714
rect 4214 82118 4266 82170
rect 4278 82118 4330 82170
rect 4342 82118 4394 82170
rect 4406 82118 4458 82170
rect 4470 82118 4522 82170
rect 34934 82118 34986 82170
rect 34998 82118 35050 82170
rect 35062 82118 35114 82170
rect 35126 82118 35178 82170
rect 35190 82118 35242 82170
rect 65654 82118 65706 82170
rect 65718 82118 65770 82170
rect 65782 82118 65834 82170
rect 65846 82118 65898 82170
rect 65910 82118 65962 82170
rect 96374 82118 96426 82170
rect 96438 82118 96490 82170
rect 96502 82118 96554 82170
rect 96566 82118 96618 82170
rect 96630 82118 96682 82170
rect 4874 81574 4926 81626
rect 4938 81574 4990 81626
rect 5002 81574 5054 81626
rect 5066 81574 5118 81626
rect 5130 81574 5182 81626
rect 35594 81574 35646 81626
rect 35658 81574 35710 81626
rect 35722 81574 35774 81626
rect 35786 81574 35838 81626
rect 35850 81574 35902 81626
rect 66314 81574 66366 81626
rect 66378 81574 66430 81626
rect 66442 81574 66494 81626
rect 66506 81574 66558 81626
rect 66570 81574 66622 81626
rect 97034 81574 97086 81626
rect 97098 81574 97150 81626
rect 97162 81574 97214 81626
rect 97226 81574 97278 81626
rect 97290 81574 97342 81626
rect 4214 81030 4266 81082
rect 4278 81030 4330 81082
rect 4342 81030 4394 81082
rect 4406 81030 4458 81082
rect 4470 81030 4522 81082
rect 34934 81030 34986 81082
rect 34998 81030 35050 81082
rect 35062 81030 35114 81082
rect 35126 81030 35178 81082
rect 35190 81030 35242 81082
rect 65654 81030 65706 81082
rect 65718 81030 65770 81082
rect 65782 81030 65834 81082
rect 65846 81030 65898 81082
rect 65910 81030 65962 81082
rect 96374 81030 96426 81082
rect 96438 81030 96490 81082
rect 96502 81030 96554 81082
rect 96566 81030 96618 81082
rect 96630 81030 96682 81082
rect 4874 80486 4926 80538
rect 4938 80486 4990 80538
rect 5002 80486 5054 80538
rect 5066 80486 5118 80538
rect 5130 80486 5182 80538
rect 35594 80486 35646 80538
rect 35658 80486 35710 80538
rect 35722 80486 35774 80538
rect 35786 80486 35838 80538
rect 35850 80486 35902 80538
rect 66314 80486 66366 80538
rect 66378 80486 66430 80538
rect 66442 80486 66494 80538
rect 66506 80486 66558 80538
rect 66570 80486 66622 80538
rect 97034 80486 97086 80538
rect 97098 80486 97150 80538
rect 97162 80486 97214 80538
rect 97226 80486 97278 80538
rect 97290 80486 97342 80538
rect 4214 79942 4266 79994
rect 4278 79942 4330 79994
rect 4342 79942 4394 79994
rect 4406 79942 4458 79994
rect 4470 79942 4522 79994
rect 34934 79942 34986 79994
rect 34998 79942 35050 79994
rect 35062 79942 35114 79994
rect 35126 79942 35178 79994
rect 35190 79942 35242 79994
rect 65654 79942 65706 79994
rect 65718 79942 65770 79994
rect 65782 79942 65834 79994
rect 65846 79942 65898 79994
rect 65910 79942 65962 79994
rect 96374 79942 96426 79994
rect 96438 79942 96490 79994
rect 96502 79942 96554 79994
rect 96566 79942 96618 79994
rect 96630 79942 96682 79994
rect 4874 79398 4926 79450
rect 4938 79398 4990 79450
rect 5002 79398 5054 79450
rect 5066 79398 5118 79450
rect 5130 79398 5182 79450
rect 35594 79398 35646 79450
rect 35658 79398 35710 79450
rect 35722 79398 35774 79450
rect 35786 79398 35838 79450
rect 35850 79398 35902 79450
rect 66314 79398 66366 79450
rect 66378 79398 66430 79450
rect 66442 79398 66494 79450
rect 66506 79398 66558 79450
rect 66570 79398 66622 79450
rect 97034 79398 97086 79450
rect 97098 79398 97150 79450
rect 97162 79398 97214 79450
rect 97226 79398 97278 79450
rect 97290 79398 97342 79450
rect 4214 78854 4266 78906
rect 4278 78854 4330 78906
rect 4342 78854 4394 78906
rect 4406 78854 4458 78906
rect 4470 78854 4522 78906
rect 34934 78854 34986 78906
rect 34998 78854 35050 78906
rect 35062 78854 35114 78906
rect 35126 78854 35178 78906
rect 35190 78854 35242 78906
rect 65654 78854 65706 78906
rect 65718 78854 65770 78906
rect 65782 78854 65834 78906
rect 65846 78854 65898 78906
rect 65910 78854 65962 78906
rect 96374 78854 96426 78906
rect 96438 78854 96490 78906
rect 96502 78854 96554 78906
rect 96566 78854 96618 78906
rect 96630 78854 96682 78906
rect 4874 78310 4926 78362
rect 4938 78310 4990 78362
rect 5002 78310 5054 78362
rect 5066 78310 5118 78362
rect 5130 78310 5182 78362
rect 35594 78310 35646 78362
rect 35658 78310 35710 78362
rect 35722 78310 35774 78362
rect 35786 78310 35838 78362
rect 35850 78310 35902 78362
rect 66314 78310 66366 78362
rect 66378 78310 66430 78362
rect 66442 78310 66494 78362
rect 66506 78310 66558 78362
rect 66570 78310 66622 78362
rect 97034 78310 97086 78362
rect 97098 78310 97150 78362
rect 97162 78310 97214 78362
rect 97226 78310 97278 78362
rect 97290 78310 97342 78362
rect 4214 77766 4266 77818
rect 4278 77766 4330 77818
rect 4342 77766 4394 77818
rect 4406 77766 4458 77818
rect 4470 77766 4522 77818
rect 34934 77766 34986 77818
rect 34998 77766 35050 77818
rect 35062 77766 35114 77818
rect 35126 77766 35178 77818
rect 35190 77766 35242 77818
rect 65654 77766 65706 77818
rect 65718 77766 65770 77818
rect 65782 77766 65834 77818
rect 65846 77766 65898 77818
rect 65910 77766 65962 77818
rect 96374 77766 96426 77818
rect 96438 77766 96490 77818
rect 96502 77766 96554 77818
rect 96566 77766 96618 77818
rect 96630 77766 96682 77818
rect 43536 77707 43588 77716
rect 43536 77673 43545 77707
rect 43545 77673 43579 77707
rect 43579 77673 43588 77707
rect 43536 77664 43588 77673
rect 47492 77707 47544 77716
rect 47492 77673 47501 77707
rect 47501 77673 47535 77707
rect 47535 77673 47544 77707
rect 47492 77664 47544 77673
rect 49700 77707 49752 77716
rect 49700 77673 49709 77707
rect 49709 77673 49743 77707
rect 49743 77673 49752 77707
rect 49700 77664 49752 77673
rect 53104 77707 53156 77716
rect 53104 77673 53113 77707
rect 53113 77673 53147 77707
rect 53147 77673 53156 77707
rect 53104 77664 53156 77673
rect 55128 77707 55180 77716
rect 55128 77673 55137 77707
rect 55137 77673 55171 77707
rect 55171 77673 55180 77707
rect 55128 77664 55180 77673
rect 57336 77707 57388 77716
rect 57336 77673 57345 77707
rect 57345 77673 57379 77707
rect 57379 77673 57388 77707
rect 57336 77664 57388 77673
rect 59176 77707 59228 77716
rect 59176 77673 59185 77707
rect 59185 77673 59219 77707
rect 59219 77673 59228 77707
rect 59176 77664 59228 77673
rect 43628 77528 43680 77580
rect 49424 77528 49476 77580
rect 41788 77324 41840 77376
rect 45652 77392 45704 77444
rect 45744 77392 45796 77444
rect 47952 77392 48004 77444
rect 51080 77392 51132 77444
rect 51264 77392 51316 77444
rect 53380 77392 53432 77444
rect 49976 77324 50028 77376
rect 53288 77324 53340 77376
rect 55588 77392 55640 77444
rect 57428 77392 57480 77444
rect 59268 77392 59320 77444
rect 56876 77324 56928 77376
rect 57520 77324 57572 77376
rect 4874 77222 4926 77274
rect 4938 77222 4990 77274
rect 5002 77222 5054 77274
rect 5066 77222 5118 77274
rect 5130 77222 5182 77274
rect 35594 77222 35646 77274
rect 35658 77222 35710 77274
rect 35722 77222 35774 77274
rect 35786 77222 35838 77274
rect 35850 77222 35902 77274
rect 66314 77222 66366 77274
rect 66378 77222 66430 77274
rect 66442 77222 66494 77274
rect 66506 77222 66558 77274
rect 66570 77222 66622 77274
rect 97034 77222 97086 77274
rect 97098 77222 97150 77274
rect 97162 77222 97214 77274
rect 97226 77222 97278 77274
rect 97290 77222 97342 77274
rect 45376 77163 45428 77172
rect 45376 77129 45385 77163
rect 45385 77129 45419 77163
rect 45419 77129 45428 77163
rect 45376 77120 45428 77129
rect 51172 77163 51224 77172
rect 51172 77129 51181 77163
rect 51181 77129 51215 77163
rect 51215 77129 51224 77163
rect 51172 77120 51224 77129
rect 48228 77052 48280 77104
rect 49608 77052 49660 77104
rect 53196 77052 53248 77104
rect 43628 77027 43680 77036
rect 43628 76993 43637 77027
rect 43637 76993 43671 77027
rect 43671 76993 43680 77027
rect 43628 76984 43680 76993
rect 49424 77027 49476 77036
rect 49424 76993 49433 77027
rect 49433 76993 49467 77027
rect 49467 76993 49476 77027
rect 49424 76984 49476 76993
rect 43628 76848 43680 76900
rect 41788 76823 41840 76832
rect 41788 76789 41797 76823
rect 41797 76789 41831 76823
rect 41831 76789 41840 76823
rect 41788 76780 41840 76789
rect 45744 76823 45796 76832
rect 45744 76789 45753 76823
rect 45753 76789 45787 76823
rect 45787 76789 45796 76823
rect 45744 76780 45796 76789
rect 47952 76823 48004 76832
rect 47952 76789 47961 76823
rect 47961 76789 47995 76823
rect 47995 76789 48004 76823
rect 47952 76780 48004 76789
rect 51264 76780 51316 76832
rect 53288 76780 53340 76832
rect 55588 76823 55640 76832
rect 55588 76789 55597 76823
rect 55597 76789 55631 76823
rect 55631 76789 55640 76823
rect 55588 76780 55640 76789
rect 57520 76823 57572 76832
rect 57520 76789 57529 76823
rect 57529 76789 57563 76823
rect 57563 76789 57572 76823
rect 57520 76780 57572 76789
rect 4214 76678 4266 76730
rect 4278 76678 4330 76730
rect 4342 76678 4394 76730
rect 4406 76678 4458 76730
rect 4470 76678 4522 76730
rect 34934 76678 34986 76730
rect 34998 76678 35050 76730
rect 35062 76678 35114 76730
rect 35126 76678 35178 76730
rect 35190 76678 35242 76730
rect 65654 76678 65706 76730
rect 65718 76678 65770 76730
rect 65782 76678 65834 76730
rect 65846 76678 65898 76730
rect 65910 76678 65962 76730
rect 96374 76678 96426 76730
rect 96438 76678 96490 76730
rect 96502 76678 96554 76730
rect 96566 76678 96618 76730
rect 96630 76678 96682 76730
rect 49608 76576 49660 76628
rect 43628 76279 43680 76288
rect 43628 76245 43637 76279
rect 43637 76245 43671 76279
rect 43671 76245 43680 76279
rect 43628 76236 43680 76245
rect 4874 76134 4926 76186
rect 4938 76134 4990 76186
rect 5002 76134 5054 76186
rect 5066 76134 5118 76186
rect 5130 76134 5182 76186
rect 35594 76134 35646 76186
rect 35658 76134 35710 76186
rect 35722 76134 35774 76186
rect 35786 76134 35838 76186
rect 35850 76134 35902 76186
rect 66314 76134 66366 76186
rect 66378 76134 66430 76186
rect 66442 76134 66494 76186
rect 66506 76134 66558 76186
rect 66570 76134 66622 76186
rect 97034 76134 97086 76186
rect 97098 76134 97150 76186
rect 97162 76134 97214 76186
rect 97226 76134 97278 76186
rect 97290 76134 97342 76186
rect 4214 75590 4266 75642
rect 4278 75590 4330 75642
rect 4342 75590 4394 75642
rect 4406 75590 4458 75642
rect 4470 75590 4522 75642
rect 34934 75590 34986 75642
rect 34998 75590 35050 75642
rect 35062 75590 35114 75642
rect 35126 75590 35178 75642
rect 35190 75590 35242 75642
rect 65654 75590 65706 75642
rect 65718 75590 65770 75642
rect 65782 75590 65834 75642
rect 65846 75590 65898 75642
rect 65910 75590 65962 75642
rect 96374 75590 96426 75642
rect 96438 75590 96490 75642
rect 96502 75590 96554 75642
rect 96566 75590 96618 75642
rect 96630 75590 96682 75642
rect 4874 75046 4926 75098
rect 4938 75046 4990 75098
rect 5002 75046 5054 75098
rect 5066 75046 5118 75098
rect 5130 75046 5182 75098
rect 35594 75046 35646 75098
rect 35658 75046 35710 75098
rect 35722 75046 35774 75098
rect 35786 75046 35838 75098
rect 35850 75046 35902 75098
rect 66314 75046 66366 75098
rect 66378 75046 66430 75098
rect 66442 75046 66494 75098
rect 66506 75046 66558 75098
rect 66570 75046 66622 75098
rect 97034 75046 97086 75098
rect 97098 75046 97150 75098
rect 97162 75046 97214 75098
rect 97226 75046 97278 75098
rect 97290 75046 97342 75098
rect 45652 74944 45704 74996
rect 48228 74987 48280 74996
rect 48228 74953 48237 74987
rect 48237 74953 48271 74987
rect 48271 74953 48280 74987
rect 48228 74944 48280 74953
rect 49976 74987 50028 74996
rect 49976 74953 49985 74987
rect 49985 74953 50019 74987
rect 50019 74953 50028 74987
rect 49976 74944 50028 74953
rect 51080 74944 51132 74996
rect 53196 74987 53248 74996
rect 53196 74953 53205 74987
rect 53205 74953 53239 74987
rect 53239 74953 53248 74987
rect 53196 74944 53248 74953
rect 53380 74944 53432 74996
rect 56876 74987 56928 74996
rect 56876 74953 56885 74987
rect 56885 74953 56919 74987
rect 56919 74953 56928 74987
rect 56876 74944 56928 74953
rect 57428 74944 57480 74996
rect 59268 74944 59320 74996
rect 46664 74851 46716 74860
rect 46664 74817 46673 74851
rect 46673 74817 46707 74851
rect 46707 74817 46716 74851
rect 46664 74808 46716 74817
rect 83924 74808 83976 74860
rect 4214 74502 4266 74554
rect 4278 74502 4330 74554
rect 4342 74502 4394 74554
rect 4406 74502 4458 74554
rect 4470 74502 4522 74554
rect 34934 74502 34986 74554
rect 34998 74502 35050 74554
rect 35062 74502 35114 74554
rect 35126 74502 35178 74554
rect 35190 74502 35242 74554
rect 65654 74502 65706 74554
rect 65718 74502 65770 74554
rect 65782 74502 65834 74554
rect 65846 74502 65898 74554
rect 65910 74502 65962 74554
rect 96374 74502 96426 74554
rect 96438 74502 96490 74554
rect 96502 74502 96554 74554
rect 96566 74502 96618 74554
rect 96630 74502 96682 74554
rect 4874 73958 4926 74010
rect 4938 73958 4990 74010
rect 5002 73958 5054 74010
rect 5066 73958 5118 74010
rect 5130 73958 5182 74010
rect 35594 73958 35646 74010
rect 35658 73958 35710 74010
rect 35722 73958 35774 74010
rect 35786 73958 35838 74010
rect 35850 73958 35902 74010
rect 66314 73958 66366 74010
rect 66378 73958 66430 74010
rect 66442 73958 66494 74010
rect 66506 73958 66558 74010
rect 66570 73958 66622 74010
rect 97034 73958 97086 74010
rect 97098 73958 97150 74010
rect 97162 73958 97214 74010
rect 97226 73958 97278 74010
rect 97290 73958 97342 74010
rect 4214 73414 4266 73466
rect 4278 73414 4330 73466
rect 4342 73414 4394 73466
rect 4406 73414 4458 73466
rect 4470 73414 4522 73466
rect 34934 73414 34986 73466
rect 34998 73414 35050 73466
rect 35062 73414 35114 73466
rect 35126 73414 35178 73466
rect 35190 73414 35242 73466
rect 65654 73414 65706 73466
rect 65718 73414 65770 73466
rect 65782 73414 65834 73466
rect 65846 73414 65898 73466
rect 65910 73414 65962 73466
rect 96374 73414 96426 73466
rect 96438 73414 96490 73466
rect 96502 73414 96554 73466
rect 96566 73414 96618 73466
rect 96630 73414 96682 73466
rect 4874 72870 4926 72922
rect 4938 72870 4990 72922
rect 5002 72870 5054 72922
rect 5066 72870 5118 72922
rect 5130 72870 5182 72922
rect 35594 72870 35646 72922
rect 35658 72870 35710 72922
rect 35722 72870 35774 72922
rect 35786 72870 35838 72922
rect 35850 72870 35902 72922
rect 66314 72870 66366 72922
rect 66378 72870 66430 72922
rect 66442 72870 66494 72922
rect 66506 72870 66558 72922
rect 66570 72870 66622 72922
rect 97034 72870 97086 72922
rect 97098 72870 97150 72922
rect 97162 72870 97214 72922
rect 97226 72870 97278 72922
rect 97290 72870 97342 72922
rect 4214 72326 4266 72378
rect 4278 72326 4330 72378
rect 4342 72326 4394 72378
rect 4406 72326 4458 72378
rect 4470 72326 4522 72378
rect 34934 72326 34986 72378
rect 34998 72326 35050 72378
rect 35062 72326 35114 72378
rect 35126 72326 35178 72378
rect 35190 72326 35242 72378
rect 65654 72326 65706 72378
rect 65718 72326 65770 72378
rect 65782 72326 65834 72378
rect 65846 72326 65898 72378
rect 65910 72326 65962 72378
rect 96374 72326 96426 72378
rect 96438 72326 96490 72378
rect 96502 72326 96554 72378
rect 96566 72326 96618 72378
rect 96630 72326 96682 72378
rect 4874 71782 4926 71834
rect 4938 71782 4990 71834
rect 5002 71782 5054 71834
rect 5066 71782 5118 71834
rect 5130 71782 5182 71834
rect 35594 71782 35646 71834
rect 35658 71782 35710 71834
rect 35722 71782 35774 71834
rect 35786 71782 35838 71834
rect 35850 71782 35902 71834
rect 66314 71782 66366 71834
rect 66378 71782 66430 71834
rect 66442 71782 66494 71834
rect 66506 71782 66558 71834
rect 66570 71782 66622 71834
rect 97034 71782 97086 71834
rect 97098 71782 97150 71834
rect 97162 71782 97214 71834
rect 97226 71782 97278 71834
rect 97290 71782 97342 71834
rect 4214 71238 4266 71290
rect 4278 71238 4330 71290
rect 4342 71238 4394 71290
rect 4406 71238 4458 71290
rect 4470 71238 4522 71290
rect 34934 71238 34986 71290
rect 34998 71238 35050 71290
rect 35062 71238 35114 71290
rect 35126 71238 35178 71290
rect 35190 71238 35242 71290
rect 65654 71238 65706 71290
rect 65718 71238 65770 71290
rect 65782 71238 65834 71290
rect 65846 71238 65898 71290
rect 65910 71238 65962 71290
rect 96374 71238 96426 71290
rect 96438 71238 96490 71290
rect 96502 71238 96554 71290
rect 96566 71238 96618 71290
rect 96630 71238 96682 71290
rect 4874 70694 4926 70746
rect 4938 70694 4990 70746
rect 5002 70694 5054 70746
rect 5066 70694 5118 70746
rect 5130 70694 5182 70746
rect 35594 70694 35646 70746
rect 35658 70694 35710 70746
rect 35722 70694 35774 70746
rect 35786 70694 35838 70746
rect 35850 70694 35902 70746
rect 66314 70694 66366 70746
rect 66378 70694 66430 70746
rect 66442 70694 66494 70746
rect 66506 70694 66558 70746
rect 66570 70694 66622 70746
rect 97034 70694 97086 70746
rect 97098 70694 97150 70746
rect 97162 70694 97214 70746
rect 97226 70694 97278 70746
rect 97290 70694 97342 70746
rect 4214 70150 4266 70202
rect 4278 70150 4330 70202
rect 4342 70150 4394 70202
rect 4406 70150 4458 70202
rect 4470 70150 4522 70202
rect 34934 70150 34986 70202
rect 34998 70150 35050 70202
rect 35062 70150 35114 70202
rect 35126 70150 35178 70202
rect 35190 70150 35242 70202
rect 65654 70150 65706 70202
rect 65718 70150 65770 70202
rect 65782 70150 65834 70202
rect 65846 70150 65898 70202
rect 65910 70150 65962 70202
rect 96374 70150 96426 70202
rect 96438 70150 96490 70202
rect 96502 70150 96554 70202
rect 96566 70150 96618 70202
rect 96630 70150 96682 70202
rect 4874 69606 4926 69658
rect 4938 69606 4990 69658
rect 5002 69606 5054 69658
rect 5066 69606 5118 69658
rect 5130 69606 5182 69658
rect 35594 69606 35646 69658
rect 35658 69606 35710 69658
rect 35722 69606 35774 69658
rect 35786 69606 35838 69658
rect 35850 69606 35902 69658
rect 66314 69606 66366 69658
rect 66378 69606 66430 69658
rect 66442 69606 66494 69658
rect 66506 69606 66558 69658
rect 66570 69606 66622 69658
rect 97034 69606 97086 69658
rect 97098 69606 97150 69658
rect 97162 69606 97214 69658
rect 97226 69606 97278 69658
rect 97290 69606 97342 69658
rect 4214 69062 4266 69114
rect 4278 69062 4330 69114
rect 4342 69062 4394 69114
rect 4406 69062 4458 69114
rect 4470 69062 4522 69114
rect 34934 69062 34986 69114
rect 34998 69062 35050 69114
rect 35062 69062 35114 69114
rect 35126 69062 35178 69114
rect 35190 69062 35242 69114
rect 65654 69062 65706 69114
rect 65718 69062 65770 69114
rect 65782 69062 65834 69114
rect 65846 69062 65898 69114
rect 65910 69062 65962 69114
rect 96374 69062 96426 69114
rect 96438 69062 96490 69114
rect 96502 69062 96554 69114
rect 96566 69062 96618 69114
rect 96630 69062 96682 69114
rect 4874 68518 4926 68570
rect 4938 68518 4990 68570
rect 5002 68518 5054 68570
rect 5066 68518 5118 68570
rect 5130 68518 5182 68570
rect 35594 68518 35646 68570
rect 35658 68518 35710 68570
rect 35722 68518 35774 68570
rect 35786 68518 35838 68570
rect 35850 68518 35902 68570
rect 66314 68518 66366 68570
rect 66378 68518 66430 68570
rect 66442 68518 66494 68570
rect 66506 68518 66558 68570
rect 66570 68518 66622 68570
rect 97034 68518 97086 68570
rect 97098 68518 97150 68570
rect 97162 68518 97214 68570
rect 97226 68518 97278 68570
rect 97290 68518 97342 68570
rect 4214 67974 4266 68026
rect 4278 67974 4330 68026
rect 4342 67974 4394 68026
rect 4406 67974 4458 68026
rect 4470 67974 4522 68026
rect 34934 67974 34986 68026
rect 34998 67974 35050 68026
rect 35062 67974 35114 68026
rect 35126 67974 35178 68026
rect 35190 67974 35242 68026
rect 65654 67974 65706 68026
rect 65718 67974 65770 68026
rect 65782 67974 65834 68026
rect 65846 67974 65898 68026
rect 65910 67974 65962 68026
rect 96374 67974 96426 68026
rect 96438 67974 96490 68026
rect 96502 67974 96554 68026
rect 96566 67974 96618 68026
rect 96630 67974 96682 68026
rect 4874 67430 4926 67482
rect 4938 67430 4990 67482
rect 5002 67430 5054 67482
rect 5066 67430 5118 67482
rect 5130 67430 5182 67482
rect 35594 67430 35646 67482
rect 35658 67430 35710 67482
rect 35722 67430 35774 67482
rect 35786 67430 35838 67482
rect 35850 67430 35902 67482
rect 66314 67430 66366 67482
rect 66378 67430 66430 67482
rect 66442 67430 66494 67482
rect 66506 67430 66558 67482
rect 66570 67430 66622 67482
rect 97034 67430 97086 67482
rect 97098 67430 97150 67482
rect 97162 67430 97214 67482
rect 97226 67430 97278 67482
rect 97290 67430 97342 67482
rect 4214 66886 4266 66938
rect 4278 66886 4330 66938
rect 4342 66886 4394 66938
rect 4406 66886 4458 66938
rect 4470 66886 4522 66938
rect 34934 66886 34986 66938
rect 34998 66886 35050 66938
rect 35062 66886 35114 66938
rect 35126 66886 35178 66938
rect 35190 66886 35242 66938
rect 65654 66886 65706 66938
rect 65718 66886 65770 66938
rect 65782 66886 65834 66938
rect 65846 66886 65898 66938
rect 65910 66886 65962 66938
rect 96374 66886 96426 66938
rect 96438 66886 96490 66938
rect 96502 66886 96554 66938
rect 96566 66886 96618 66938
rect 96630 66886 96682 66938
rect 4874 66342 4926 66394
rect 4938 66342 4990 66394
rect 5002 66342 5054 66394
rect 5066 66342 5118 66394
rect 5130 66342 5182 66394
rect 35594 66342 35646 66394
rect 35658 66342 35710 66394
rect 35722 66342 35774 66394
rect 35786 66342 35838 66394
rect 35850 66342 35902 66394
rect 66314 66342 66366 66394
rect 66378 66342 66430 66394
rect 66442 66342 66494 66394
rect 66506 66342 66558 66394
rect 66570 66342 66622 66394
rect 97034 66342 97086 66394
rect 97098 66342 97150 66394
rect 97162 66342 97214 66394
rect 97226 66342 97278 66394
rect 97290 66342 97342 66394
rect 4214 65798 4266 65850
rect 4278 65798 4330 65850
rect 4342 65798 4394 65850
rect 4406 65798 4458 65850
rect 4470 65798 4522 65850
rect 34934 65798 34986 65850
rect 34998 65798 35050 65850
rect 35062 65798 35114 65850
rect 35126 65798 35178 65850
rect 35190 65798 35242 65850
rect 65654 65798 65706 65850
rect 65718 65798 65770 65850
rect 65782 65798 65834 65850
rect 65846 65798 65898 65850
rect 65910 65798 65962 65850
rect 96374 65798 96426 65850
rect 96438 65798 96490 65850
rect 96502 65798 96554 65850
rect 96566 65798 96618 65850
rect 96630 65798 96682 65850
rect 4874 65254 4926 65306
rect 4938 65254 4990 65306
rect 5002 65254 5054 65306
rect 5066 65254 5118 65306
rect 5130 65254 5182 65306
rect 35594 65254 35646 65306
rect 35658 65254 35710 65306
rect 35722 65254 35774 65306
rect 35786 65254 35838 65306
rect 35850 65254 35902 65306
rect 66314 65254 66366 65306
rect 66378 65254 66430 65306
rect 66442 65254 66494 65306
rect 66506 65254 66558 65306
rect 66570 65254 66622 65306
rect 97034 65254 97086 65306
rect 97098 65254 97150 65306
rect 97162 65254 97214 65306
rect 97226 65254 97278 65306
rect 97290 65254 97342 65306
rect 4214 64710 4266 64762
rect 4278 64710 4330 64762
rect 4342 64710 4394 64762
rect 4406 64710 4458 64762
rect 4470 64710 4522 64762
rect 34934 64710 34986 64762
rect 34998 64710 35050 64762
rect 35062 64710 35114 64762
rect 35126 64710 35178 64762
rect 35190 64710 35242 64762
rect 65654 64710 65706 64762
rect 65718 64710 65770 64762
rect 65782 64710 65834 64762
rect 65846 64710 65898 64762
rect 65910 64710 65962 64762
rect 96374 64710 96426 64762
rect 96438 64710 96490 64762
rect 96502 64710 96554 64762
rect 96566 64710 96618 64762
rect 96630 64710 96682 64762
rect 4874 64166 4926 64218
rect 4938 64166 4990 64218
rect 5002 64166 5054 64218
rect 5066 64166 5118 64218
rect 5130 64166 5182 64218
rect 35594 64166 35646 64218
rect 35658 64166 35710 64218
rect 35722 64166 35774 64218
rect 35786 64166 35838 64218
rect 35850 64166 35902 64218
rect 66314 64166 66366 64218
rect 66378 64166 66430 64218
rect 66442 64166 66494 64218
rect 66506 64166 66558 64218
rect 66570 64166 66622 64218
rect 97034 64166 97086 64218
rect 97098 64166 97150 64218
rect 97162 64166 97214 64218
rect 97226 64166 97278 64218
rect 97290 64166 97342 64218
rect 4214 63622 4266 63674
rect 4278 63622 4330 63674
rect 4342 63622 4394 63674
rect 4406 63622 4458 63674
rect 4470 63622 4522 63674
rect 34934 63622 34986 63674
rect 34998 63622 35050 63674
rect 35062 63622 35114 63674
rect 35126 63622 35178 63674
rect 35190 63622 35242 63674
rect 65654 63622 65706 63674
rect 65718 63622 65770 63674
rect 65782 63622 65834 63674
rect 65846 63622 65898 63674
rect 65910 63622 65962 63674
rect 96374 63622 96426 63674
rect 96438 63622 96490 63674
rect 96502 63622 96554 63674
rect 96566 63622 96618 63674
rect 96630 63622 96682 63674
rect 4874 63078 4926 63130
rect 4938 63078 4990 63130
rect 5002 63078 5054 63130
rect 5066 63078 5118 63130
rect 5130 63078 5182 63130
rect 35594 63078 35646 63130
rect 35658 63078 35710 63130
rect 35722 63078 35774 63130
rect 35786 63078 35838 63130
rect 35850 63078 35902 63130
rect 66314 63078 66366 63130
rect 66378 63078 66430 63130
rect 66442 63078 66494 63130
rect 66506 63078 66558 63130
rect 66570 63078 66622 63130
rect 97034 63078 97086 63130
rect 97098 63078 97150 63130
rect 97162 63078 97214 63130
rect 97226 63078 97278 63130
rect 97290 63078 97342 63130
rect 96252 62840 96304 62892
rect 100392 62679 100444 62688
rect 100392 62645 100401 62679
rect 100401 62645 100435 62679
rect 100435 62645 100444 62679
rect 100392 62636 100444 62645
rect 4214 62534 4266 62586
rect 4278 62534 4330 62586
rect 4342 62534 4394 62586
rect 4406 62534 4458 62586
rect 4470 62534 4522 62586
rect 34934 62534 34986 62586
rect 34998 62534 35050 62586
rect 35062 62534 35114 62586
rect 35126 62534 35178 62586
rect 35190 62534 35242 62586
rect 65654 62534 65706 62586
rect 65718 62534 65770 62586
rect 65782 62534 65834 62586
rect 65846 62534 65898 62586
rect 65910 62534 65962 62586
rect 96374 62534 96426 62586
rect 96438 62534 96490 62586
rect 96502 62534 96554 62586
rect 96566 62534 96618 62586
rect 96630 62534 96682 62586
rect 96896 62228 96948 62280
rect 1492 62135 1544 62144
rect 1492 62101 1501 62135
rect 1501 62101 1535 62135
rect 1535 62101 1544 62135
rect 1492 62092 1544 62101
rect 1860 62135 1912 62144
rect 1860 62101 1869 62135
rect 1869 62101 1903 62135
rect 1903 62101 1912 62135
rect 1860 62092 1912 62101
rect 100392 62135 100444 62144
rect 100392 62101 100401 62135
rect 100401 62101 100435 62135
rect 100435 62101 100444 62135
rect 100392 62092 100444 62101
rect 4874 61990 4926 62042
rect 4938 61990 4990 62042
rect 5002 61990 5054 62042
rect 5066 61990 5118 62042
rect 5130 61990 5182 62042
rect 35594 61990 35646 62042
rect 35658 61990 35710 62042
rect 35722 61990 35774 62042
rect 35786 61990 35838 62042
rect 35850 61990 35902 62042
rect 66314 61990 66366 62042
rect 66378 61990 66430 62042
rect 66442 61990 66494 62042
rect 66506 61990 66558 62042
rect 66570 61990 66622 62042
rect 97034 61990 97086 62042
rect 97098 61990 97150 62042
rect 97162 61990 97214 62042
rect 97226 61990 97278 62042
rect 97290 61990 97342 62042
rect 21088 61752 21140 61804
rect 100208 61795 100260 61804
rect 100208 61761 100217 61795
rect 100217 61761 100251 61795
rect 100251 61761 100260 61795
rect 100208 61752 100260 61761
rect 848 61548 900 61600
rect 100392 61591 100444 61600
rect 100392 61557 100401 61591
rect 100401 61557 100435 61591
rect 100435 61557 100444 61591
rect 100392 61548 100444 61557
rect 4214 61446 4266 61498
rect 4278 61446 4330 61498
rect 4342 61446 4394 61498
rect 4406 61446 4458 61498
rect 4470 61446 4522 61498
rect 34934 61446 34986 61498
rect 34998 61446 35050 61498
rect 35062 61446 35114 61498
rect 35126 61446 35178 61498
rect 35190 61446 35242 61498
rect 65654 61446 65706 61498
rect 65718 61446 65770 61498
rect 65782 61446 65834 61498
rect 65846 61446 65898 61498
rect 65910 61446 65962 61498
rect 96374 61446 96426 61498
rect 96438 61446 96490 61498
rect 96502 61446 96554 61498
rect 96566 61446 96618 61498
rect 96630 61446 96682 61498
rect 21088 61387 21140 61396
rect 21088 61353 21097 61387
rect 21097 61353 21131 61387
rect 21131 61353 21140 61387
rect 21088 61344 21140 61353
rect 77116 61344 77168 61396
rect 82452 61344 82504 61396
rect 96252 61344 96304 61396
rect 28172 61208 28224 61260
rect 79692 61208 79744 61260
rect 79876 61208 79928 61260
rect 22836 61183 22888 61192
rect 22836 61149 22845 61183
rect 22845 61149 22879 61183
rect 22879 61149 22888 61183
rect 22836 61140 22888 61149
rect 77024 61183 77076 61192
rect 77024 61149 77033 61183
rect 77033 61149 77067 61183
rect 77067 61149 77076 61183
rect 77024 61140 77076 61149
rect 96896 61208 96948 61260
rect 81532 61140 81584 61192
rect 83924 61183 83976 61192
rect 83924 61149 83933 61183
rect 83933 61149 83967 61183
rect 83967 61149 83976 61183
rect 83924 61140 83976 61149
rect 28816 61004 28868 61056
rect 71780 61004 71832 61056
rect 77760 61072 77812 61124
rect 79140 61115 79192 61124
rect 79140 61081 79149 61115
rect 79149 61081 79183 61115
rect 79183 61081 79192 61115
rect 79140 61072 79192 61081
rect 79600 61072 79652 61124
rect 82452 61072 82504 61124
rect 82820 61072 82872 61124
rect 83832 61047 83884 61056
rect 83832 61013 83841 61047
rect 83841 61013 83875 61047
rect 83875 61013 83884 61047
rect 83832 61004 83884 61013
rect 84016 61047 84068 61056
rect 84016 61013 84025 61047
rect 84025 61013 84059 61047
rect 84059 61013 84068 61047
rect 84016 61004 84068 61013
rect 4874 60902 4926 60954
rect 4938 60902 4990 60954
rect 5002 60902 5054 60954
rect 5066 60902 5118 60954
rect 5130 60902 5182 60954
rect 35594 60902 35646 60954
rect 35658 60902 35710 60954
rect 35722 60902 35774 60954
rect 35786 60902 35838 60954
rect 35850 60902 35902 60954
rect 66314 60902 66366 60954
rect 66378 60902 66430 60954
rect 66442 60902 66494 60954
rect 66506 60902 66558 60954
rect 66570 60902 66622 60954
rect 97034 60902 97086 60954
rect 97098 60902 97150 60954
rect 97162 60902 97214 60954
rect 97226 60902 97278 60954
rect 97290 60902 97342 60954
rect 79140 60800 79192 60852
rect 79876 60800 79928 60852
rect 83832 60800 83884 60852
rect 24032 60639 24084 60648
rect 24032 60605 24041 60639
rect 24041 60605 24075 60639
rect 24075 60605 24084 60639
rect 24032 60596 24084 60605
rect 48412 60732 48464 60784
rect 49424 60732 49476 60784
rect 28816 60664 28868 60716
rect 46664 60664 46716 60716
rect 79232 60707 79284 60716
rect 79232 60673 79241 60707
rect 79241 60673 79275 60707
rect 79275 60673 79284 60707
rect 79232 60664 79284 60673
rect 81716 60732 81768 60784
rect 84016 60732 84068 60784
rect 85580 60732 85632 60784
rect 79692 60707 79744 60716
rect 79692 60673 79701 60707
rect 79701 60673 79735 60707
rect 79735 60673 79744 60707
rect 79692 60664 79744 60673
rect 1860 60460 1912 60512
rect 22376 60503 22428 60512
rect 22376 60469 22385 60503
rect 22385 60469 22419 60503
rect 22419 60469 22428 60503
rect 22376 60460 22428 60469
rect 22836 60460 22888 60512
rect 77760 60596 77812 60648
rect 79600 60596 79652 60648
rect 81532 60639 81584 60648
rect 81532 60605 81541 60639
rect 81541 60605 81575 60639
rect 81575 60605 81584 60639
rect 81532 60596 81584 60605
rect 81808 60639 81860 60648
rect 81808 60605 81817 60639
rect 81817 60605 81851 60639
rect 81851 60605 81860 60639
rect 81808 60596 81860 60605
rect 83924 60639 83976 60648
rect 83924 60605 83933 60639
rect 83933 60605 83967 60639
rect 83967 60605 83976 60639
rect 83924 60596 83976 60605
rect 85672 60639 85724 60648
rect 85672 60605 85681 60639
rect 85681 60605 85715 60639
rect 85715 60605 85724 60639
rect 85672 60596 85724 60605
rect 79508 60503 79560 60512
rect 79508 60469 79517 60503
rect 79517 60469 79551 60503
rect 79551 60469 79560 60503
rect 79508 60460 79560 60469
rect 79692 60460 79744 60512
rect 81440 60503 81492 60512
rect 81440 60469 81449 60503
rect 81449 60469 81483 60503
rect 81483 60469 81492 60503
rect 81440 60460 81492 60469
rect 83280 60503 83332 60512
rect 83280 60469 83289 60503
rect 83289 60469 83323 60503
rect 83323 60469 83332 60503
rect 83280 60460 83332 60469
rect 86132 60503 86184 60512
rect 86132 60469 86141 60503
rect 86141 60469 86175 60503
rect 86175 60469 86184 60503
rect 86132 60460 86184 60469
rect 87604 60639 87656 60648
rect 87604 60605 87613 60639
rect 87613 60605 87647 60639
rect 87647 60605 87656 60639
rect 87604 60596 87656 60605
rect 87880 60639 87932 60648
rect 87880 60605 87889 60639
rect 87889 60605 87923 60639
rect 87923 60605 87932 60639
rect 87880 60596 87932 60605
rect 100392 60571 100444 60580
rect 100392 60537 100401 60571
rect 100401 60537 100435 60571
rect 100435 60537 100444 60571
rect 100392 60528 100444 60537
rect 87880 60460 87932 60512
rect 1322 60358 1374 60410
rect 1386 60358 1438 60410
rect 4214 60358 4266 60410
rect 4278 60358 4330 60410
rect 4342 60358 4394 60410
rect 4406 60358 4458 60410
rect 4470 60358 4522 60410
rect 34934 60358 34986 60410
rect 34998 60358 35050 60410
rect 35062 60358 35114 60410
rect 35126 60358 35178 60410
rect 35190 60358 35242 60410
rect 65654 60358 65706 60410
rect 65718 60358 65770 60410
rect 65782 60358 65834 60410
rect 65846 60358 65898 60410
rect 65910 60358 65962 60410
rect 96374 60358 96426 60410
rect 96438 60358 96490 60410
rect 96502 60358 96554 60410
rect 96566 60358 96618 60410
rect 96630 60358 96682 60410
rect 98930 60358 98982 60410
rect 98994 60358 99046 60410
rect 99058 60358 99110 60410
rect 99122 60358 99174 60410
rect 99186 60358 99238 60410
rect 24032 60256 24084 60308
rect 29184 60256 29236 60308
rect 48412 60299 48464 60308
rect 48412 60265 48421 60299
rect 48421 60265 48455 60299
rect 48455 60265 48464 60299
rect 48412 60256 48464 60265
rect 81716 60256 81768 60308
rect 82820 60256 82872 60308
rect 85580 60256 85632 60308
rect 85672 60256 85724 60308
rect 87604 60256 87656 60308
rect 83280 60188 83332 60240
rect 100208 60256 100260 60308
rect 91744 60188 91796 60240
rect 77024 60120 77076 60172
rect 83924 60120 83976 60172
rect 79232 60052 79284 60104
rect 81348 60052 81400 60104
rect 83832 60052 83884 60104
rect 84384 60095 84436 60104
rect 84384 60061 84393 60095
rect 84393 60061 84427 60095
rect 84427 60061 84436 60095
rect 84384 60052 84436 60061
rect 86132 60052 86184 60104
rect 89536 60052 89588 60104
rect 89720 60052 89772 60104
rect 98368 60052 98420 60104
rect 57060 60027 57112 60036
rect 57060 59993 57069 60027
rect 57069 59993 57103 60027
rect 57103 59993 57112 60027
rect 57060 59984 57112 59993
rect 81440 59984 81492 60036
rect 91744 59984 91796 60036
rect 100392 59959 100444 59968
rect 100392 59925 100401 59959
rect 100401 59925 100435 59959
rect 100435 59925 100444 59959
rect 100392 59916 100444 59925
rect 1690 59814 1742 59866
rect 1754 59814 1806 59866
rect 4874 59814 4926 59866
rect 4938 59814 4990 59866
rect 5002 59814 5054 59866
rect 5066 59814 5118 59866
rect 5130 59814 5182 59866
rect 35594 59814 35646 59866
rect 35658 59814 35710 59866
rect 35722 59814 35774 59866
rect 35786 59814 35838 59866
rect 35850 59814 35902 59866
rect 66314 59814 66366 59866
rect 66378 59814 66430 59866
rect 66442 59814 66494 59866
rect 66506 59814 66558 59866
rect 66570 59814 66622 59866
rect 97034 59814 97086 59866
rect 97098 59814 97150 59866
rect 97162 59814 97214 59866
rect 97226 59814 97278 59866
rect 97290 59814 97342 59866
rect 99666 59814 99718 59866
rect 99730 59814 99782 59866
rect 99794 59814 99846 59866
rect 99858 59814 99910 59866
rect 99922 59814 99974 59866
rect 2688 59372 2740 59424
rect 22376 59372 22428 59424
rect 1322 59270 1374 59322
rect 1386 59270 1438 59322
rect 98930 59270 98982 59322
rect 98994 59270 99046 59322
rect 99058 59270 99110 59322
rect 99122 59270 99174 59322
rect 99186 59270 99238 59322
rect 1690 58726 1742 58778
rect 1754 58726 1806 58778
rect 84384 58760 84436 58812
rect 97356 58760 97408 58812
rect 81348 58692 81400 58744
rect 97448 58692 97500 58744
rect 99666 58726 99718 58778
rect 99730 58726 99782 58778
rect 99794 58726 99846 58778
rect 99858 58726 99910 58778
rect 99922 58726 99974 58778
rect 57060 58624 57112 58676
rect 97264 58624 97316 58676
rect 1322 58182 1374 58234
rect 1386 58182 1438 58234
rect 98930 58182 98982 58234
rect 98994 58182 99046 58234
rect 99058 58182 99110 58234
rect 99122 58182 99174 58234
rect 99186 58182 99238 58234
rect 1690 57638 1742 57690
rect 1754 57638 1806 57690
rect 99666 57638 99718 57690
rect 99730 57638 99782 57690
rect 99794 57638 99846 57690
rect 99858 57638 99910 57690
rect 99922 57638 99974 57690
rect 1322 57094 1374 57146
rect 1386 57094 1438 57146
rect 98930 57094 98982 57146
rect 98994 57094 99046 57146
rect 99058 57094 99110 57146
rect 99122 57094 99174 57146
rect 99186 57094 99238 57146
rect 1690 56550 1742 56602
rect 1754 56550 1806 56602
rect 99666 56550 99718 56602
rect 99730 56550 99782 56602
rect 99794 56550 99846 56602
rect 99858 56550 99910 56602
rect 99922 56550 99974 56602
rect 1322 56006 1374 56058
rect 1386 56006 1438 56058
rect 98930 56006 98982 56058
rect 98994 56006 99046 56058
rect 99058 56006 99110 56058
rect 99122 56006 99174 56058
rect 99186 56006 99238 56058
rect 1690 55462 1742 55514
rect 1754 55462 1806 55514
rect 99666 55462 99718 55514
rect 99730 55462 99782 55514
rect 99794 55462 99846 55514
rect 99858 55462 99910 55514
rect 99922 55462 99974 55514
rect 1322 54918 1374 54970
rect 1386 54918 1438 54970
rect 98930 54918 98982 54970
rect 98994 54918 99046 54970
rect 99058 54918 99110 54970
rect 99122 54918 99174 54970
rect 99186 54918 99238 54970
rect 1690 54374 1742 54426
rect 1754 54374 1806 54426
rect 99666 54374 99718 54426
rect 99730 54374 99782 54426
rect 99794 54374 99846 54426
rect 99858 54374 99910 54426
rect 99922 54374 99974 54426
rect 97080 53932 97132 53984
rect 1322 53830 1374 53882
rect 1386 53830 1438 53882
rect 98930 53830 98982 53882
rect 98994 53830 99046 53882
rect 99058 53830 99110 53882
rect 99122 53830 99174 53882
rect 99186 53830 99238 53882
rect 1690 53286 1742 53338
rect 1754 53286 1806 53338
rect 99666 53286 99718 53338
rect 99730 53286 99782 53338
rect 99794 53286 99846 53338
rect 99858 53286 99910 53338
rect 99922 53286 99974 53338
rect 1322 52742 1374 52794
rect 1386 52742 1438 52794
rect 98930 52742 98982 52794
rect 98994 52742 99046 52794
rect 99058 52742 99110 52794
rect 99122 52742 99174 52794
rect 99186 52742 99238 52794
rect 1690 52198 1742 52250
rect 1754 52198 1806 52250
rect 99666 52198 99718 52250
rect 99730 52198 99782 52250
rect 99794 52198 99846 52250
rect 99858 52198 99910 52250
rect 99922 52198 99974 52250
rect 1322 51654 1374 51706
rect 1386 51654 1438 51706
rect 98930 51654 98982 51706
rect 98994 51654 99046 51706
rect 99058 51654 99110 51706
rect 99122 51654 99174 51706
rect 99186 51654 99238 51706
rect 1690 51110 1742 51162
rect 1754 51110 1806 51162
rect 99666 51110 99718 51162
rect 99730 51110 99782 51162
rect 99794 51110 99846 51162
rect 99858 51110 99910 51162
rect 99922 51110 99974 51162
rect 1322 50566 1374 50618
rect 1386 50566 1438 50618
rect 98930 50566 98982 50618
rect 98994 50566 99046 50618
rect 99058 50566 99110 50618
rect 99122 50566 99174 50618
rect 99186 50566 99238 50618
rect 1690 50022 1742 50074
rect 1754 50022 1806 50074
rect 99666 50022 99718 50074
rect 99730 50022 99782 50074
rect 99794 50022 99846 50074
rect 99858 50022 99910 50074
rect 99922 50022 99974 50074
rect 1322 49478 1374 49530
rect 1386 49478 1438 49530
rect 98930 49478 98982 49530
rect 98994 49478 99046 49530
rect 99058 49478 99110 49530
rect 99122 49478 99174 49530
rect 99186 49478 99238 49530
rect 1690 48934 1742 48986
rect 1754 48934 1806 48986
rect 99666 48934 99718 48986
rect 99730 48934 99782 48986
rect 99794 48934 99846 48986
rect 99858 48934 99910 48986
rect 99922 48934 99974 48986
rect 1322 48390 1374 48442
rect 1386 48390 1438 48442
rect 98930 48390 98982 48442
rect 98994 48390 99046 48442
rect 99058 48390 99110 48442
rect 99122 48390 99174 48442
rect 99186 48390 99238 48442
rect 1690 47846 1742 47898
rect 1754 47846 1806 47898
rect 99666 47846 99718 47898
rect 99730 47846 99782 47898
rect 99794 47846 99846 47898
rect 99858 47846 99910 47898
rect 99922 47846 99974 47898
rect 1322 47302 1374 47354
rect 1386 47302 1438 47354
rect 98930 47302 98982 47354
rect 98994 47302 99046 47354
rect 99058 47302 99110 47354
rect 99122 47302 99174 47354
rect 99186 47302 99238 47354
rect 1690 46758 1742 46810
rect 1754 46758 1806 46810
rect 99666 46758 99718 46810
rect 99730 46758 99782 46810
rect 99794 46758 99846 46810
rect 99858 46758 99910 46810
rect 99922 46758 99974 46810
rect 1322 46214 1374 46266
rect 1386 46214 1438 46266
rect 98930 46214 98982 46266
rect 98994 46214 99046 46266
rect 99058 46214 99110 46266
rect 99122 46214 99174 46266
rect 99186 46214 99238 46266
rect 98552 46087 98604 46096
rect 98552 46053 98561 46087
rect 98561 46053 98595 46087
rect 98595 46053 98604 46087
rect 98552 46044 98604 46053
rect 98276 45951 98328 45960
rect 98276 45917 98285 45951
rect 98285 45917 98319 45951
rect 98319 45917 98328 45951
rect 98276 45908 98328 45917
rect 98368 45951 98420 45960
rect 98368 45917 98377 45951
rect 98377 45917 98411 45951
rect 98411 45917 98420 45951
rect 98368 45908 98420 45917
rect 98184 45840 98236 45892
rect 1690 45670 1742 45722
rect 1754 45670 1806 45722
rect 99666 45670 99718 45722
rect 99730 45670 99782 45722
rect 99794 45670 99846 45722
rect 99858 45670 99910 45722
rect 99922 45670 99974 45722
rect 1322 45126 1374 45178
rect 1386 45126 1438 45178
rect 98930 45126 98982 45178
rect 98994 45126 99046 45178
rect 99058 45126 99110 45178
rect 99122 45126 99174 45178
rect 99186 45126 99238 45178
rect 98276 45024 98328 45076
rect 98368 44752 98420 44804
rect 98184 44684 98236 44736
rect 98644 44727 98696 44736
rect 98644 44693 98653 44727
rect 98653 44693 98687 44727
rect 98687 44693 98696 44727
rect 98644 44684 98696 44693
rect 1690 44582 1742 44634
rect 1754 44582 1806 44634
rect 99666 44582 99718 44634
rect 99730 44582 99782 44634
rect 99794 44582 99846 44634
rect 99858 44582 99910 44634
rect 99922 44582 99974 44634
rect 1322 44038 1374 44090
rect 1386 44038 1438 44090
rect 98930 44038 98982 44090
rect 98994 44038 99046 44090
rect 99058 44038 99110 44090
rect 99122 44038 99174 44090
rect 99186 44038 99238 44090
rect 1690 43494 1742 43546
rect 1754 43494 1806 43546
rect 99666 43494 99718 43546
rect 99730 43494 99782 43546
rect 99794 43494 99846 43546
rect 99858 43494 99910 43546
rect 99922 43494 99974 43546
rect 97448 43256 97500 43308
rect 98276 43299 98328 43308
rect 98276 43265 98285 43299
rect 98285 43265 98319 43299
rect 98319 43265 98328 43299
rect 98276 43256 98328 43265
rect 98368 43095 98420 43104
rect 98368 43061 98377 43095
rect 98377 43061 98411 43095
rect 98411 43061 98420 43095
rect 98368 43052 98420 43061
rect 1322 42950 1374 43002
rect 1386 42950 1438 43002
rect 98930 42950 98982 43002
rect 98994 42950 99046 43002
rect 99058 42950 99110 43002
rect 99122 42950 99174 43002
rect 99186 42950 99238 43002
rect 1690 42406 1742 42458
rect 1754 42406 1806 42458
rect 99666 42406 99718 42458
rect 99730 42406 99782 42458
rect 99794 42406 99846 42458
rect 99858 42406 99910 42458
rect 99922 42406 99974 42458
rect 1322 41862 1374 41914
rect 1386 41862 1438 41914
rect 98930 41862 98982 41914
rect 98994 41862 99046 41914
rect 99058 41862 99110 41914
rect 99122 41862 99174 41914
rect 99186 41862 99238 41914
rect 1690 41318 1742 41370
rect 1754 41318 1806 41370
rect 99666 41318 99718 41370
rect 99730 41318 99782 41370
rect 99794 41318 99846 41370
rect 99858 41318 99910 41370
rect 99922 41318 99974 41370
rect 98368 41148 98420 41200
rect 98460 41012 98512 41064
rect 100116 41055 100168 41064
rect 100116 41021 100125 41055
rect 100125 41021 100159 41055
rect 100159 41021 100168 41055
rect 100116 41012 100168 41021
rect 98184 40876 98236 40928
rect 1322 40774 1374 40826
rect 1386 40774 1438 40826
rect 98930 40774 98982 40826
rect 98994 40774 99046 40826
rect 99058 40774 99110 40826
rect 99122 40774 99174 40826
rect 99186 40774 99238 40826
rect 98460 40715 98512 40724
rect 98460 40681 98469 40715
rect 98469 40681 98503 40715
rect 98503 40681 98512 40715
rect 98460 40672 98512 40681
rect 98552 40468 98604 40520
rect 98644 40400 98696 40452
rect 100208 40400 100260 40452
rect 1690 40230 1742 40282
rect 1754 40230 1806 40282
rect 99666 40230 99718 40282
rect 99730 40230 99782 40282
rect 99794 40230 99846 40282
rect 99858 40230 99910 40282
rect 99922 40230 99974 40282
rect 1322 39686 1374 39738
rect 1386 39686 1438 39738
rect 98930 39686 98982 39738
rect 98994 39686 99046 39738
rect 99058 39686 99110 39738
rect 99122 39686 99174 39738
rect 99186 39686 99238 39738
rect 1690 39142 1742 39194
rect 1754 39142 1806 39194
rect 99666 39142 99718 39194
rect 99730 39142 99782 39194
rect 99794 39142 99846 39194
rect 99858 39142 99910 39194
rect 99922 39142 99974 39194
rect 1322 38598 1374 38650
rect 1386 38598 1438 38650
rect 98930 38598 98982 38650
rect 98994 38598 99046 38650
rect 99058 38598 99110 38650
rect 99122 38598 99174 38650
rect 99186 38598 99238 38650
rect 1690 38054 1742 38106
rect 1754 38054 1806 38106
rect 99666 38054 99718 38106
rect 99730 38054 99782 38106
rect 99794 38054 99846 38106
rect 99858 38054 99910 38106
rect 99922 38054 99974 38106
rect 1322 37510 1374 37562
rect 1386 37510 1438 37562
rect 98930 37510 98982 37562
rect 98994 37510 99046 37562
rect 99058 37510 99110 37562
rect 99122 37510 99174 37562
rect 99186 37510 99238 37562
rect 1690 36966 1742 37018
rect 1754 36966 1806 37018
rect 99666 36966 99718 37018
rect 99730 36966 99782 37018
rect 99794 36966 99846 37018
rect 99858 36966 99910 37018
rect 99922 36966 99974 37018
rect 1322 36422 1374 36474
rect 1386 36422 1438 36474
rect 98930 36422 98982 36474
rect 98994 36422 99046 36474
rect 99058 36422 99110 36474
rect 99122 36422 99174 36474
rect 99186 36422 99238 36474
rect 1690 35878 1742 35930
rect 1754 35878 1806 35930
rect 99666 35878 99718 35930
rect 99730 35878 99782 35930
rect 99794 35878 99846 35930
rect 99858 35878 99910 35930
rect 99922 35878 99974 35930
rect 98276 35683 98328 35692
rect 98276 35649 98285 35683
rect 98285 35649 98319 35683
rect 98319 35649 98328 35683
rect 98276 35640 98328 35649
rect 98460 35640 98512 35692
rect 98736 35436 98788 35488
rect 1322 35334 1374 35386
rect 1386 35334 1438 35386
rect 98930 35334 98982 35386
rect 98994 35334 99046 35386
rect 99058 35334 99110 35386
rect 99122 35334 99174 35386
rect 99186 35334 99238 35386
rect 1690 34790 1742 34842
rect 1754 34790 1806 34842
rect 99666 34790 99718 34842
rect 99730 34790 99782 34842
rect 99794 34790 99846 34842
rect 99858 34790 99910 34842
rect 99922 34790 99974 34842
rect 98460 34552 98512 34604
rect 98368 34527 98420 34536
rect 98368 34493 98377 34527
rect 98377 34493 98411 34527
rect 98411 34493 98420 34527
rect 98368 34484 98420 34493
rect 1322 34246 1374 34298
rect 1386 34246 1438 34298
rect 98930 34246 98982 34298
rect 98994 34246 99046 34298
rect 99058 34246 99110 34298
rect 99122 34246 99174 34298
rect 99186 34246 99238 34298
rect 1690 33702 1742 33754
rect 1754 33702 1806 33754
rect 99666 33702 99718 33754
rect 99730 33702 99782 33754
rect 99794 33702 99846 33754
rect 99858 33702 99910 33754
rect 99922 33702 99974 33754
rect 1322 33158 1374 33210
rect 1386 33158 1438 33210
rect 98930 33158 98982 33210
rect 98994 33158 99046 33210
rect 99058 33158 99110 33210
rect 99122 33158 99174 33210
rect 99186 33158 99238 33210
rect 1690 32614 1742 32666
rect 1754 32614 1806 32666
rect 99666 32614 99718 32666
rect 99730 32614 99782 32666
rect 99794 32614 99846 32666
rect 99858 32614 99910 32666
rect 99922 32614 99974 32666
rect 1322 32070 1374 32122
rect 1386 32070 1438 32122
rect 98930 32070 98982 32122
rect 98994 32070 99046 32122
rect 99058 32070 99110 32122
rect 99122 32070 99174 32122
rect 99186 32070 99238 32122
rect 99380 31832 99432 31884
rect 99840 31875 99892 31884
rect 99840 31841 99849 31875
rect 99849 31841 99883 31875
rect 99883 31841 99892 31875
rect 99840 31832 99892 31841
rect 98736 31764 98788 31816
rect 100208 31764 100260 31816
rect 1690 31526 1742 31578
rect 1754 31526 1806 31578
rect 99666 31526 99718 31578
rect 99730 31526 99782 31578
rect 99794 31526 99846 31578
rect 99858 31526 99910 31578
rect 99922 31526 99974 31578
rect 1322 30982 1374 31034
rect 1386 30982 1438 31034
rect 98930 30982 98982 31034
rect 98994 30982 99046 31034
rect 99058 30982 99110 31034
rect 99122 30982 99174 31034
rect 99186 30982 99238 31034
rect 100208 30676 100260 30728
rect 98368 30608 98420 30660
rect 98276 30583 98328 30592
rect 98276 30549 98285 30583
rect 98285 30549 98319 30583
rect 98319 30549 98328 30583
rect 98276 30540 98328 30549
rect 99564 30540 99616 30592
rect 1690 30438 1742 30490
rect 1754 30438 1806 30490
rect 99666 30438 99718 30490
rect 99730 30438 99782 30490
rect 99794 30438 99846 30490
rect 99858 30438 99910 30490
rect 99922 30438 99974 30490
rect 99380 30200 99432 30252
rect 100116 30200 100168 30252
rect 99380 30039 99432 30048
rect 99380 30005 99389 30039
rect 99389 30005 99423 30039
rect 99423 30005 99432 30039
rect 99380 29996 99432 30005
rect 1322 29894 1374 29946
rect 1386 29894 1438 29946
rect 98930 29894 98982 29946
rect 98994 29894 99046 29946
rect 99058 29894 99110 29946
rect 99122 29894 99174 29946
rect 99186 29894 99238 29946
rect 98460 29588 98512 29640
rect 98736 29588 98788 29640
rect 98644 29452 98696 29504
rect 1690 29350 1742 29402
rect 1754 29350 1806 29402
rect 99666 29350 99718 29402
rect 99730 29350 99782 29402
rect 99794 29350 99846 29402
rect 99858 29350 99910 29402
rect 99922 29350 99974 29402
rect 98736 29112 98788 29164
rect 99380 29112 99432 29164
rect 98276 29044 98328 29096
rect 99288 29044 99340 29096
rect 100300 29044 100352 29096
rect 98552 28976 98604 29028
rect 99472 29019 99524 29028
rect 99472 28985 99481 29019
rect 99481 28985 99515 29019
rect 99515 28985 99524 29019
rect 99472 28976 99524 28985
rect 100024 28976 100076 29028
rect 1322 28806 1374 28858
rect 1386 28806 1438 28858
rect 98930 28806 98982 28858
rect 98994 28806 99046 28858
rect 99058 28806 99110 28858
rect 99122 28806 99174 28858
rect 99186 28806 99238 28858
rect 1690 28262 1742 28314
rect 1754 28262 1806 28314
rect 99666 28262 99718 28314
rect 99730 28262 99782 28314
rect 99794 28262 99846 28314
rect 99858 28262 99910 28314
rect 99922 28262 99974 28314
rect 1322 27718 1374 27770
rect 1386 27718 1438 27770
rect 98930 27718 98982 27770
rect 98994 27718 99046 27770
rect 99058 27718 99110 27770
rect 99122 27718 99174 27770
rect 99186 27718 99238 27770
rect 97356 27548 97408 27600
rect 98368 27548 98420 27600
rect 99564 27548 99616 27600
rect 99472 27412 99524 27464
rect 99564 27344 99616 27396
rect 100024 27412 100076 27464
rect 100300 27412 100352 27464
rect 100116 27344 100168 27396
rect 1690 27174 1742 27226
rect 1754 27174 1806 27226
rect 99666 27174 99718 27226
rect 99730 27174 99782 27226
rect 99794 27174 99846 27226
rect 99858 27174 99910 27226
rect 99922 27174 99974 27226
rect 1322 26630 1374 26682
rect 1386 26630 1438 26682
rect 98930 26630 98982 26682
rect 98994 26630 99046 26682
rect 99058 26630 99110 26682
rect 99122 26630 99174 26682
rect 99186 26630 99238 26682
rect 98368 26392 98420 26444
rect 100484 26367 100536 26376
rect 100484 26333 100493 26367
rect 100493 26333 100527 26367
rect 100527 26333 100536 26367
rect 100484 26324 100536 26333
rect 1690 26086 1742 26138
rect 1754 26086 1806 26138
rect 99666 26086 99718 26138
rect 99730 26086 99782 26138
rect 99794 26086 99846 26138
rect 99858 26086 99910 26138
rect 99922 26086 99974 26138
rect 100024 25984 100076 26036
rect 98368 25959 98420 25968
rect 98368 25925 98377 25959
rect 98377 25925 98411 25959
rect 98411 25925 98420 25959
rect 98368 25916 98420 25925
rect 99564 25848 99616 25900
rect 98368 25780 98420 25832
rect 98736 25780 98788 25832
rect 98828 25712 98880 25764
rect 99288 25712 99340 25764
rect 98276 25644 98328 25696
rect 1322 25542 1374 25594
rect 1386 25542 1438 25594
rect 98930 25542 98982 25594
rect 98994 25542 99046 25594
rect 99058 25542 99110 25594
rect 99122 25542 99174 25594
rect 99186 25542 99238 25594
rect 98644 25304 98696 25356
rect 99288 25304 99340 25356
rect 100208 25236 100260 25288
rect 98092 25100 98144 25152
rect 1690 24998 1742 25050
rect 1754 24998 1806 25050
rect 99666 24998 99718 25050
rect 99730 24998 99782 25050
rect 99794 24998 99846 25050
rect 99858 24998 99910 25050
rect 99922 24998 99974 25050
rect 98552 24760 98604 24812
rect 99380 24692 99432 24744
rect 100208 24735 100260 24744
rect 100208 24701 100217 24735
rect 100217 24701 100251 24735
rect 100251 24701 100260 24735
rect 100208 24692 100260 24701
rect 98552 24556 98604 24608
rect 1322 24454 1374 24506
rect 1386 24454 1438 24506
rect 98930 24454 98982 24506
rect 98994 24454 99046 24506
rect 99058 24454 99110 24506
rect 99122 24454 99174 24506
rect 99186 24454 99238 24506
rect 98368 24191 98420 24200
rect 98368 24157 98377 24191
rect 98377 24157 98411 24191
rect 98411 24157 98420 24191
rect 98368 24148 98420 24157
rect 98460 24055 98512 24064
rect 98460 24021 98469 24055
rect 98469 24021 98503 24055
rect 98503 24021 98512 24055
rect 98460 24012 98512 24021
rect 1690 23910 1742 23962
rect 1754 23910 1806 23962
rect 99666 23910 99718 23962
rect 99730 23910 99782 23962
rect 99794 23910 99846 23962
rect 99858 23910 99910 23962
rect 99922 23910 99974 23962
rect 98736 23851 98788 23860
rect 98736 23817 98745 23851
rect 98745 23817 98779 23851
rect 98779 23817 98788 23851
rect 98736 23808 98788 23817
rect 99288 23808 99340 23860
rect 98276 23715 98328 23724
rect 98276 23681 98285 23715
rect 98285 23681 98319 23715
rect 98319 23681 98328 23715
rect 98276 23672 98328 23681
rect 99472 23672 99524 23724
rect 100024 23672 100076 23724
rect 98092 23468 98144 23520
rect 98368 23511 98420 23520
rect 98368 23477 98377 23511
rect 98377 23477 98411 23511
rect 98411 23477 98420 23511
rect 98368 23468 98420 23477
rect 1322 23366 1374 23418
rect 1386 23366 1438 23418
rect 98930 23366 98982 23418
rect 98994 23366 99046 23418
rect 99058 23366 99110 23418
rect 99122 23366 99174 23418
rect 99186 23366 99238 23418
rect 1690 22822 1742 22874
rect 1754 22822 1806 22874
rect 99666 22822 99718 22874
rect 99730 22822 99782 22874
rect 99794 22822 99846 22874
rect 99858 22822 99910 22874
rect 99922 22822 99974 22874
rect 97356 22720 97408 22772
rect 98368 22720 98420 22772
rect 98736 22720 98788 22772
rect 99380 22763 99432 22772
rect 99380 22729 99389 22763
rect 99389 22729 99423 22763
rect 99423 22729 99432 22763
rect 99380 22720 99432 22729
rect 99472 22720 99524 22772
rect 98276 22516 98328 22568
rect 98552 22516 98604 22568
rect 99288 22627 99340 22636
rect 99288 22593 99297 22627
rect 99297 22593 99331 22627
rect 99331 22593 99340 22627
rect 99288 22584 99340 22593
rect 98552 22380 98604 22432
rect 98828 22380 98880 22432
rect 99380 22380 99432 22432
rect 99564 22380 99616 22432
rect 1322 22278 1374 22330
rect 1386 22278 1438 22330
rect 98930 22278 98982 22330
rect 98994 22278 99046 22330
rect 99058 22278 99110 22330
rect 99122 22278 99174 22330
rect 99186 22278 99238 22330
rect 99472 22176 99524 22228
rect 97540 21904 97592 21956
rect 98276 21947 98328 21956
rect 98276 21913 98285 21947
rect 98285 21913 98319 21947
rect 98319 21913 98328 21947
rect 98276 21904 98328 21913
rect 98736 21904 98788 21956
rect 98644 21879 98696 21888
rect 98644 21845 98653 21879
rect 98653 21845 98687 21879
rect 98687 21845 98696 21879
rect 98644 21836 98696 21845
rect 99288 21836 99340 21888
rect 1690 21734 1742 21786
rect 1754 21734 1806 21786
rect 99666 21734 99718 21786
rect 99730 21734 99782 21786
rect 99794 21734 99846 21786
rect 99858 21734 99910 21786
rect 99922 21734 99974 21786
rect 1322 21190 1374 21242
rect 1386 21190 1438 21242
rect 98930 21190 98982 21242
rect 98994 21190 99046 21242
rect 99058 21190 99110 21242
rect 99122 21190 99174 21242
rect 99186 21190 99238 21242
rect 1690 20646 1742 20698
rect 1754 20646 1806 20698
rect 99666 20646 99718 20698
rect 99730 20646 99782 20698
rect 99794 20646 99846 20698
rect 99858 20646 99910 20698
rect 99922 20646 99974 20698
rect 1322 20102 1374 20154
rect 1386 20102 1438 20154
rect 98930 20102 98982 20154
rect 98994 20102 99046 20154
rect 99058 20102 99110 20154
rect 99122 20102 99174 20154
rect 99186 20102 99238 20154
rect 98828 19864 98880 19916
rect 100208 19864 100260 19916
rect 98460 19728 98512 19780
rect 98368 19703 98420 19712
rect 98368 19669 98377 19703
rect 98377 19669 98411 19703
rect 98411 19669 98420 19703
rect 98368 19660 98420 19669
rect 1690 19558 1742 19610
rect 1754 19558 1806 19610
rect 99666 19558 99718 19610
rect 99730 19558 99782 19610
rect 99794 19558 99846 19610
rect 99858 19558 99910 19610
rect 99922 19558 99974 19610
rect 98368 19252 98420 19304
rect 98460 19159 98512 19168
rect 98460 19125 98469 19159
rect 98469 19125 98503 19159
rect 98503 19125 98512 19159
rect 98460 19116 98512 19125
rect 1322 19014 1374 19066
rect 1386 19014 1438 19066
rect 98930 19014 98982 19066
rect 98994 19014 99046 19066
rect 99058 19014 99110 19066
rect 99122 19014 99174 19066
rect 99186 19014 99238 19066
rect 1690 18470 1742 18522
rect 1754 18470 1806 18522
rect 99666 18470 99718 18522
rect 99730 18470 99782 18522
rect 99794 18470 99846 18522
rect 99858 18470 99910 18522
rect 99922 18470 99974 18522
rect 98460 18275 98512 18284
rect 98460 18241 98469 18275
rect 98469 18241 98503 18275
rect 98503 18241 98512 18275
rect 98460 18232 98512 18241
rect 98644 18164 98696 18216
rect 98828 18207 98880 18216
rect 98828 18173 98837 18207
rect 98837 18173 98871 18207
rect 98871 18173 98880 18207
rect 98828 18164 98880 18173
rect 1322 17926 1374 17978
rect 1386 17926 1438 17978
rect 98930 17926 98982 17978
rect 98994 17926 99046 17978
rect 99058 17926 99110 17978
rect 99122 17926 99174 17978
rect 99186 17926 99238 17978
rect 1690 17382 1742 17434
rect 1754 17382 1806 17434
rect 99666 17382 99718 17434
rect 99730 17382 99782 17434
rect 99794 17382 99846 17434
rect 99858 17382 99910 17434
rect 99922 17382 99974 17434
rect 1322 16838 1374 16890
rect 1386 16838 1438 16890
rect 98930 16838 98982 16890
rect 98994 16838 99046 16890
rect 99058 16838 99110 16890
rect 99122 16838 99174 16890
rect 99186 16838 99238 16890
rect 1690 16294 1742 16346
rect 1754 16294 1806 16346
rect 99666 16294 99718 16346
rect 99730 16294 99782 16346
rect 99794 16294 99846 16346
rect 99858 16294 99910 16346
rect 99922 16294 99974 16346
rect 1322 15750 1374 15802
rect 1386 15750 1438 15802
rect 98930 15750 98982 15802
rect 98994 15750 99046 15802
rect 99058 15750 99110 15802
rect 99122 15750 99174 15802
rect 99186 15750 99238 15802
rect 1690 15206 1742 15258
rect 1754 15206 1806 15258
rect 99666 15206 99718 15258
rect 99730 15206 99782 15258
rect 99794 15206 99846 15258
rect 99858 15206 99910 15258
rect 99922 15206 99974 15258
rect 1322 14662 1374 14714
rect 1386 14662 1438 14714
rect 98930 14662 98982 14714
rect 98994 14662 99046 14714
rect 99058 14662 99110 14714
rect 99122 14662 99174 14714
rect 99186 14662 99238 14714
rect 1690 14118 1742 14170
rect 1754 14118 1806 14170
rect 99666 14118 99718 14170
rect 99730 14118 99782 14170
rect 99794 14118 99846 14170
rect 99858 14118 99910 14170
rect 99922 14118 99974 14170
rect 1322 13574 1374 13626
rect 1386 13574 1438 13626
rect 98930 13574 98982 13626
rect 98994 13574 99046 13626
rect 99058 13574 99110 13626
rect 99122 13574 99174 13626
rect 99186 13574 99238 13626
rect 1690 13030 1742 13082
rect 1754 13030 1806 13082
rect 99666 13030 99718 13082
rect 99730 13030 99782 13082
rect 99794 13030 99846 13082
rect 99858 13030 99910 13082
rect 99922 13030 99974 13082
rect 1322 12486 1374 12538
rect 1386 12486 1438 12538
rect 98930 12486 98982 12538
rect 98994 12486 99046 12538
rect 99058 12486 99110 12538
rect 99122 12486 99174 12538
rect 99186 12486 99238 12538
rect 1690 11942 1742 11994
rect 1754 11942 1806 11994
rect 99666 11942 99718 11994
rect 99730 11942 99782 11994
rect 99794 11942 99846 11994
rect 99858 11942 99910 11994
rect 99922 11942 99974 11994
rect 1322 11398 1374 11450
rect 1386 11398 1438 11450
rect 98930 11398 98982 11450
rect 98994 11398 99046 11450
rect 99058 11398 99110 11450
rect 99122 11398 99174 11450
rect 99186 11398 99238 11450
rect 1690 10854 1742 10906
rect 1754 10854 1806 10906
rect 99666 10854 99718 10906
rect 99730 10854 99782 10906
rect 99794 10854 99846 10906
rect 99858 10854 99910 10906
rect 99922 10854 99974 10906
rect 1322 10310 1374 10362
rect 1386 10310 1438 10362
rect 98930 10310 98982 10362
rect 98994 10310 99046 10362
rect 99058 10310 99110 10362
rect 99122 10310 99174 10362
rect 99186 10310 99238 10362
rect 1690 9766 1742 9818
rect 1754 9766 1806 9818
rect 99666 9766 99718 9818
rect 99730 9766 99782 9818
rect 99794 9766 99846 9818
rect 99858 9766 99910 9818
rect 99922 9766 99974 9818
rect 1322 9222 1374 9274
rect 1386 9222 1438 9274
rect 98930 9222 98982 9274
rect 98994 9222 99046 9274
rect 99058 9222 99110 9274
rect 99122 9222 99174 9274
rect 99186 9222 99238 9274
rect 1690 8678 1742 8730
rect 1754 8678 1806 8730
rect 99666 8678 99718 8730
rect 99730 8678 99782 8730
rect 99794 8678 99846 8730
rect 99858 8678 99910 8730
rect 99922 8678 99974 8730
rect 1322 8134 1374 8186
rect 1386 8134 1438 8186
rect 98930 8134 98982 8186
rect 98994 8134 99046 8186
rect 99058 8134 99110 8186
rect 99122 8134 99174 8186
rect 99186 8134 99238 8186
rect 1690 7590 1742 7642
rect 1754 7590 1806 7642
rect 99666 7590 99718 7642
rect 99730 7590 99782 7642
rect 99794 7590 99846 7642
rect 99858 7590 99910 7642
rect 99922 7590 99974 7642
rect 1322 7046 1374 7098
rect 1386 7046 1438 7098
rect 98930 7046 98982 7098
rect 98994 7046 99046 7098
rect 99058 7046 99110 7098
rect 99122 7046 99174 7098
rect 99186 7046 99238 7098
rect 1690 6502 1742 6554
rect 1754 6502 1806 6554
rect 99666 6502 99718 6554
rect 99730 6502 99782 6554
rect 99794 6502 99846 6554
rect 99858 6502 99910 6554
rect 99922 6502 99974 6554
rect 1322 5958 1374 6010
rect 1386 5958 1438 6010
rect 98930 5958 98982 6010
rect 98994 5958 99046 6010
rect 99058 5958 99110 6010
rect 99122 5958 99174 6010
rect 99186 5958 99238 6010
rect 1690 5414 1742 5466
rect 1754 5414 1806 5466
rect 99666 5414 99718 5466
rect 99730 5414 99782 5466
rect 99794 5414 99846 5466
rect 99858 5414 99910 5466
rect 99922 5414 99974 5466
rect 1322 4870 1374 4922
rect 1386 4870 1438 4922
rect 98930 4870 98982 4922
rect 98994 4870 99046 4922
rect 99058 4870 99110 4922
rect 99122 4870 99174 4922
rect 99186 4870 99238 4922
rect 1690 4326 1742 4378
rect 1754 4326 1806 4378
rect 99666 4326 99718 4378
rect 99730 4326 99782 4378
rect 99794 4326 99846 4378
rect 99858 4326 99910 4378
rect 99922 4326 99974 4378
rect 1322 3782 1374 3834
rect 1386 3782 1438 3834
rect 98930 3782 98982 3834
rect 98994 3782 99046 3834
rect 99058 3782 99110 3834
rect 99122 3782 99174 3834
rect 99186 3782 99238 3834
rect 1690 3238 1742 3290
rect 1754 3238 1806 3290
rect 99666 3238 99718 3290
rect 99730 3238 99782 3290
rect 99794 3238 99846 3290
rect 99858 3238 99910 3290
rect 99922 3238 99974 3290
rect 1322 2694 1374 2746
rect 1386 2694 1438 2746
rect 98930 2694 98982 2746
rect 98994 2694 99046 2746
rect 99058 2694 99110 2746
rect 99122 2694 99174 2746
rect 99186 2694 99238 2746
rect 1690 2150 1742 2202
rect 1754 2150 1806 2202
rect 99666 2150 99718 2202
rect 99730 2150 99782 2202
rect 99794 2150 99846 2202
rect 99858 2150 99910 2202
rect 99922 2150 99974 2202
<< metal2 >>
rect 43166 103442 43222 104106
rect 45098 103442 45154 104106
rect 47674 103442 47730 104106
rect 49606 103442 49662 104106
rect 43166 103414 43392 103442
rect 43166 103306 43222 103414
rect 4214 101756 4522 101765
rect 4214 101754 4220 101756
rect 4276 101754 4300 101756
rect 4356 101754 4380 101756
rect 4436 101754 4460 101756
rect 4516 101754 4522 101756
rect 4276 101702 4278 101754
rect 4458 101702 4460 101754
rect 4214 101700 4220 101702
rect 4276 101700 4300 101702
rect 4356 101700 4380 101702
rect 4436 101700 4460 101702
rect 4516 101700 4522 101702
rect 4214 101691 4522 101700
rect 34934 101756 35242 101765
rect 34934 101754 34940 101756
rect 34996 101754 35020 101756
rect 35076 101754 35100 101756
rect 35156 101754 35180 101756
rect 35236 101754 35242 101756
rect 34996 101702 34998 101754
rect 35178 101702 35180 101754
rect 34934 101700 34940 101702
rect 34996 101700 35020 101702
rect 35076 101700 35100 101702
rect 35156 101700 35180 101702
rect 35236 101700 35242 101702
rect 34934 101691 35242 101700
rect 43364 101658 43392 103414
rect 45098 103414 45324 103442
rect 45098 103306 45154 103414
rect 45296 101658 45324 103414
rect 47674 103414 47992 103442
rect 47674 103306 47730 103414
rect 47964 101658 47992 103414
rect 49528 103414 49662 103442
rect 49528 101658 49556 103414
rect 49606 103306 49662 103414
rect 50894 103442 50950 104106
rect 52826 103442 52882 104106
rect 55402 103442 55458 104106
rect 57334 103442 57390 104106
rect 58622 103442 58678 104106
rect 50894 103414 51028 103442
rect 50894 103306 50950 103414
rect 51000 101658 51028 103414
rect 52826 103414 53052 103442
rect 52826 103306 52882 103414
rect 53024 101658 53052 103414
rect 55402 103414 55720 103442
rect 55402 103306 55458 103414
rect 55692 101658 55720 103414
rect 57334 103414 57652 103442
rect 57334 103306 57390 103414
rect 57624 101658 57652 103414
rect 58622 103414 58848 103442
rect 58622 103306 58678 103414
rect 58820 101658 58848 103414
rect 65654 101756 65962 101765
rect 65654 101754 65660 101756
rect 65716 101754 65740 101756
rect 65796 101754 65820 101756
rect 65876 101754 65900 101756
rect 65956 101754 65962 101756
rect 65716 101702 65718 101754
rect 65898 101702 65900 101754
rect 65654 101700 65660 101702
rect 65716 101700 65740 101702
rect 65796 101700 65820 101702
rect 65876 101700 65900 101702
rect 65956 101700 65962 101702
rect 65654 101691 65962 101700
rect 96374 101756 96682 101765
rect 96374 101754 96380 101756
rect 96436 101754 96460 101756
rect 96516 101754 96540 101756
rect 96596 101754 96620 101756
rect 96676 101754 96682 101756
rect 96436 101702 96438 101754
rect 96618 101702 96620 101754
rect 96374 101700 96380 101702
rect 96436 101700 96460 101702
rect 96516 101700 96540 101702
rect 96596 101700 96620 101702
rect 96676 101700 96682 101702
rect 96374 101691 96682 101700
rect 43352 101652 43404 101658
rect 43352 101594 43404 101600
rect 45284 101652 45336 101658
rect 45284 101594 45336 101600
rect 47952 101652 48004 101658
rect 47952 101594 48004 101600
rect 49516 101652 49568 101658
rect 49516 101594 49568 101600
rect 50988 101652 51040 101658
rect 50988 101594 51040 101600
rect 53012 101652 53064 101658
rect 53012 101594 53064 101600
rect 55680 101652 55732 101658
rect 55680 101594 55732 101600
rect 57612 101652 57664 101658
rect 57612 101594 57664 101600
rect 58808 101652 58860 101658
rect 58808 101594 58860 101600
rect 43536 101448 43588 101454
rect 43536 101390 43588 101396
rect 45376 101448 45428 101454
rect 45376 101390 45428 101396
rect 47492 101448 47544 101454
rect 47492 101390 47544 101396
rect 49700 101448 49752 101454
rect 49700 101390 49752 101396
rect 51172 101448 51224 101454
rect 51172 101390 51224 101396
rect 53104 101448 53156 101454
rect 53104 101390 53156 101396
rect 55128 101448 55180 101454
rect 55128 101390 55180 101396
rect 57336 101448 57388 101454
rect 57336 101390 57388 101396
rect 59176 101448 59228 101454
rect 59176 101390 59228 101396
rect 4874 101212 5182 101221
rect 4874 101210 4880 101212
rect 4936 101210 4960 101212
rect 5016 101210 5040 101212
rect 5096 101210 5120 101212
rect 5176 101210 5182 101212
rect 4936 101158 4938 101210
rect 5118 101158 5120 101210
rect 4874 101156 4880 101158
rect 4936 101156 4960 101158
rect 5016 101156 5040 101158
rect 5096 101156 5120 101158
rect 5176 101156 5182 101158
rect 4874 101147 5182 101156
rect 35594 101212 35902 101221
rect 35594 101210 35600 101212
rect 35656 101210 35680 101212
rect 35736 101210 35760 101212
rect 35816 101210 35840 101212
rect 35896 101210 35902 101212
rect 35656 101158 35658 101210
rect 35838 101158 35840 101210
rect 35594 101156 35600 101158
rect 35656 101156 35680 101158
rect 35736 101156 35760 101158
rect 35816 101156 35840 101158
rect 35896 101156 35902 101158
rect 35594 101147 35902 101156
rect 4214 100668 4522 100677
rect 4214 100666 4220 100668
rect 4276 100666 4300 100668
rect 4356 100666 4380 100668
rect 4436 100666 4460 100668
rect 4516 100666 4522 100668
rect 4276 100614 4278 100666
rect 4458 100614 4460 100666
rect 4214 100612 4220 100614
rect 4276 100612 4300 100614
rect 4356 100612 4380 100614
rect 4436 100612 4460 100614
rect 4516 100612 4522 100614
rect 4214 100603 4522 100612
rect 34934 100668 35242 100677
rect 34934 100666 34940 100668
rect 34996 100666 35020 100668
rect 35076 100666 35100 100668
rect 35156 100666 35180 100668
rect 35236 100666 35242 100668
rect 34996 100614 34998 100666
rect 35178 100614 35180 100666
rect 34934 100612 34940 100614
rect 34996 100612 35020 100614
rect 35076 100612 35100 100614
rect 35156 100612 35180 100614
rect 35236 100612 35242 100614
rect 34934 100603 35242 100612
rect 4874 100124 5182 100133
rect 4874 100122 4880 100124
rect 4936 100122 4960 100124
rect 5016 100122 5040 100124
rect 5096 100122 5120 100124
rect 5176 100122 5182 100124
rect 4936 100070 4938 100122
rect 5118 100070 5120 100122
rect 4874 100068 4880 100070
rect 4936 100068 4960 100070
rect 5016 100068 5040 100070
rect 5096 100068 5120 100070
rect 5176 100068 5182 100070
rect 4874 100059 5182 100068
rect 35594 100124 35902 100133
rect 35594 100122 35600 100124
rect 35656 100122 35680 100124
rect 35736 100122 35760 100124
rect 35816 100122 35840 100124
rect 35896 100122 35902 100124
rect 35656 100070 35658 100122
rect 35838 100070 35840 100122
rect 35594 100068 35600 100070
rect 35656 100068 35680 100070
rect 35736 100068 35760 100070
rect 35816 100068 35840 100070
rect 35896 100068 35902 100070
rect 35594 100059 35902 100068
rect 4214 99580 4522 99589
rect 4214 99578 4220 99580
rect 4276 99578 4300 99580
rect 4356 99578 4380 99580
rect 4436 99578 4460 99580
rect 4516 99578 4522 99580
rect 4276 99526 4278 99578
rect 4458 99526 4460 99578
rect 4214 99524 4220 99526
rect 4276 99524 4300 99526
rect 4356 99524 4380 99526
rect 4436 99524 4460 99526
rect 4516 99524 4522 99526
rect 4214 99515 4522 99524
rect 34934 99580 35242 99589
rect 34934 99578 34940 99580
rect 34996 99578 35020 99580
rect 35076 99578 35100 99580
rect 35156 99578 35180 99580
rect 35236 99578 35242 99580
rect 34996 99526 34998 99578
rect 35178 99526 35180 99578
rect 34934 99524 34940 99526
rect 34996 99524 35020 99526
rect 35076 99524 35100 99526
rect 35156 99524 35180 99526
rect 35236 99524 35242 99526
rect 34934 99515 35242 99524
rect 4874 99036 5182 99045
rect 4874 99034 4880 99036
rect 4936 99034 4960 99036
rect 5016 99034 5040 99036
rect 5096 99034 5120 99036
rect 5176 99034 5182 99036
rect 4936 98982 4938 99034
rect 5118 98982 5120 99034
rect 4874 98980 4880 98982
rect 4936 98980 4960 98982
rect 5016 98980 5040 98982
rect 5096 98980 5120 98982
rect 5176 98980 5182 98982
rect 4874 98971 5182 98980
rect 35594 99036 35902 99045
rect 35594 99034 35600 99036
rect 35656 99034 35680 99036
rect 35736 99034 35760 99036
rect 35816 99034 35840 99036
rect 35896 99034 35902 99036
rect 35656 98982 35658 99034
rect 35838 98982 35840 99034
rect 35594 98980 35600 98982
rect 35656 98980 35680 98982
rect 35736 98980 35760 98982
rect 35816 98980 35840 98982
rect 35896 98980 35902 98982
rect 35594 98971 35902 98980
rect 4214 98492 4522 98501
rect 4214 98490 4220 98492
rect 4276 98490 4300 98492
rect 4356 98490 4380 98492
rect 4436 98490 4460 98492
rect 4516 98490 4522 98492
rect 4276 98438 4278 98490
rect 4458 98438 4460 98490
rect 4214 98436 4220 98438
rect 4276 98436 4300 98438
rect 4356 98436 4380 98438
rect 4436 98436 4460 98438
rect 4516 98436 4522 98438
rect 4214 98427 4522 98436
rect 34934 98492 35242 98501
rect 34934 98490 34940 98492
rect 34996 98490 35020 98492
rect 35076 98490 35100 98492
rect 35156 98490 35180 98492
rect 35236 98490 35242 98492
rect 34996 98438 34998 98490
rect 35178 98438 35180 98490
rect 34934 98436 34940 98438
rect 34996 98436 35020 98438
rect 35076 98436 35100 98438
rect 35156 98436 35180 98438
rect 35236 98436 35242 98438
rect 34934 98427 35242 98436
rect 4874 97948 5182 97957
rect 4874 97946 4880 97948
rect 4936 97946 4960 97948
rect 5016 97946 5040 97948
rect 5096 97946 5120 97948
rect 5176 97946 5182 97948
rect 4936 97894 4938 97946
rect 5118 97894 5120 97946
rect 4874 97892 4880 97894
rect 4936 97892 4960 97894
rect 5016 97892 5040 97894
rect 5096 97892 5120 97894
rect 5176 97892 5182 97894
rect 4874 97883 5182 97892
rect 35594 97948 35902 97957
rect 35594 97946 35600 97948
rect 35656 97946 35680 97948
rect 35736 97946 35760 97948
rect 35816 97946 35840 97948
rect 35896 97946 35902 97948
rect 35656 97894 35658 97946
rect 35838 97894 35840 97946
rect 35594 97892 35600 97894
rect 35656 97892 35680 97894
rect 35736 97892 35760 97894
rect 35816 97892 35840 97894
rect 35896 97892 35902 97894
rect 35594 97883 35902 97892
rect 4214 97404 4522 97413
rect 4214 97402 4220 97404
rect 4276 97402 4300 97404
rect 4356 97402 4380 97404
rect 4436 97402 4460 97404
rect 4516 97402 4522 97404
rect 4276 97350 4278 97402
rect 4458 97350 4460 97402
rect 4214 97348 4220 97350
rect 4276 97348 4300 97350
rect 4356 97348 4380 97350
rect 4436 97348 4460 97350
rect 4516 97348 4522 97350
rect 4214 97339 4522 97348
rect 34934 97404 35242 97413
rect 34934 97402 34940 97404
rect 34996 97402 35020 97404
rect 35076 97402 35100 97404
rect 35156 97402 35180 97404
rect 35236 97402 35242 97404
rect 34996 97350 34998 97402
rect 35178 97350 35180 97402
rect 34934 97348 34940 97350
rect 34996 97348 35020 97350
rect 35076 97348 35100 97350
rect 35156 97348 35180 97350
rect 35236 97348 35242 97350
rect 34934 97339 35242 97348
rect 4874 96860 5182 96869
rect 4874 96858 4880 96860
rect 4936 96858 4960 96860
rect 5016 96858 5040 96860
rect 5096 96858 5120 96860
rect 5176 96858 5182 96860
rect 4936 96806 4938 96858
rect 5118 96806 5120 96858
rect 4874 96804 4880 96806
rect 4936 96804 4960 96806
rect 5016 96804 5040 96806
rect 5096 96804 5120 96806
rect 5176 96804 5182 96806
rect 4874 96795 5182 96804
rect 35594 96860 35902 96869
rect 35594 96858 35600 96860
rect 35656 96858 35680 96860
rect 35736 96858 35760 96860
rect 35816 96858 35840 96860
rect 35896 96858 35902 96860
rect 35656 96806 35658 96858
rect 35838 96806 35840 96858
rect 35594 96804 35600 96806
rect 35656 96804 35680 96806
rect 35736 96804 35760 96806
rect 35816 96804 35840 96806
rect 35896 96804 35902 96806
rect 35594 96795 35902 96804
rect 4214 96316 4522 96325
rect 4214 96314 4220 96316
rect 4276 96314 4300 96316
rect 4356 96314 4380 96316
rect 4436 96314 4460 96316
rect 4516 96314 4522 96316
rect 4276 96262 4278 96314
rect 4458 96262 4460 96314
rect 4214 96260 4220 96262
rect 4276 96260 4300 96262
rect 4356 96260 4380 96262
rect 4436 96260 4460 96262
rect 4516 96260 4522 96262
rect 4214 96251 4522 96260
rect 34934 96316 35242 96325
rect 34934 96314 34940 96316
rect 34996 96314 35020 96316
rect 35076 96314 35100 96316
rect 35156 96314 35180 96316
rect 35236 96314 35242 96316
rect 34996 96262 34998 96314
rect 35178 96262 35180 96314
rect 34934 96260 34940 96262
rect 34996 96260 35020 96262
rect 35076 96260 35100 96262
rect 35156 96260 35180 96262
rect 35236 96260 35242 96262
rect 34934 96251 35242 96260
rect 4874 95772 5182 95781
rect 4874 95770 4880 95772
rect 4936 95770 4960 95772
rect 5016 95770 5040 95772
rect 5096 95770 5120 95772
rect 5176 95770 5182 95772
rect 4936 95718 4938 95770
rect 5118 95718 5120 95770
rect 4874 95716 4880 95718
rect 4936 95716 4960 95718
rect 5016 95716 5040 95718
rect 5096 95716 5120 95718
rect 5176 95716 5182 95718
rect 4874 95707 5182 95716
rect 35594 95772 35902 95781
rect 35594 95770 35600 95772
rect 35656 95770 35680 95772
rect 35736 95770 35760 95772
rect 35816 95770 35840 95772
rect 35896 95770 35902 95772
rect 35656 95718 35658 95770
rect 35838 95718 35840 95770
rect 35594 95716 35600 95718
rect 35656 95716 35680 95718
rect 35736 95716 35760 95718
rect 35816 95716 35840 95718
rect 35896 95716 35902 95718
rect 35594 95707 35902 95716
rect 4214 95228 4522 95237
rect 4214 95226 4220 95228
rect 4276 95226 4300 95228
rect 4356 95226 4380 95228
rect 4436 95226 4460 95228
rect 4516 95226 4522 95228
rect 4276 95174 4278 95226
rect 4458 95174 4460 95226
rect 4214 95172 4220 95174
rect 4276 95172 4300 95174
rect 4356 95172 4380 95174
rect 4436 95172 4460 95174
rect 4516 95172 4522 95174
rect 4214 95163 4522 95172
rect 34934 95228 35242 95237
rect 34934 95226 34940 95228
rect 34996 95226 35020 95228
rect 35076 95226 35100 95228
rect 35156 95226 35180 95228
rect 35236 95226 35242 95228
rect 34996 95174 34998 95226
rect 35178 95174 35180 95226
rect 34934 95172 34940 95174
rect 34996 95172 35020 95174
rect 35076 95172 35100 95174
rect 35156 95172 35180 95174
rect 35236 95172 35242 95174
rect 34934 95163 35242 95172
rect 4874 94684 5182 94693
rect 4874 94682 4880 94684
rect 4936 94682 4960 94684
rect 5016 94682 5040 94684
rect 5096 94682 5120 94684
rect 5176 94682 5182 94684
rect 4936 94630 4938 94682
rect 5118 94630 5120 94682
rect 4874 94628 4880 94630
rect 4936 94628 4960 94630
rect 5016 94628 5040 94630
rect 5096 94628 5120 94630
rect 5176 94628 5182 94630
rect 4874 94619 5182 94628
rect 35594 94684 35902 94693
rect 35594 94682 35600 94684
rect 35656 94682 35680 94684
rect 35736 94682 35760 94684
rect 35816 94682 35840 94684
rect 35896 94682 35902 94684
rect 35656 94630 35658 94682
rect 35838 94630 35840 94682
rect 35594 94628 35600 94630
rect 35656 94628 35680 94630
rect 35736 94628 35760 94630
rect 35816 94628 35840 94630
rect 35896 94628 35902 94630
rect 35594 94619 35902 94628
rect 4214 94140 4522 94149
rect 4214 94138 4220 94140
rect 4276 94138 4300 94140
rect 4356 94138 4380 94140
rect 4436 94138 4460 94140
rect 4516 94138 4522 94140
rect 4276 94086 4278 94138
rect 4458 94086 4460 94138
rect 4214 94084 4220 94086
rect 4276 94084 4300 94086
rect 4356 94084 4380 94086
rect 4436 94084 4460 94086
rect 4516 94084 4522 94086
rect 4214 94075 4522 94084
rect 34934 94140 35242 94149
rect 34934 94138 34940 94140
rect 34996 94138 35020 94140
rect 35076 94138 35100 94140
rect 35156 94138 35180 94140
rect 35236 94138 35242 94140
rect 34996 94086 34998 94138
rect 35178 94086 35180 94138
rect 34934 94084 34940 94086
rect 34996 94084 35020 94086
rect 35076 94084 35100 94086
rect 35156 94084 35180 94086
rect 35236 94084 35242 94086
rect 34934 94075 35242 94084
rect 4874 93596 5182 93605
rect 4874 93594 4880 93596
rect 4936 93594 4960 93596
rect 5016 93594 5040 93596
rect 5096 93594 5120 93596
rect 5176 93594 5182 93596
rect 4936 93542 4938 93594
rect 5118 93542 5120 93594
rect 4874 93540 4880 93542
rect 4936 93540 4960 93542
rect 5016 93540 5040 93542
rect 5096 93540 5120 93542
rect 5176 93540 5182 93542
rect 4874 93531 5182 93540
rect 35594 93596 35902 93605
rect 35594 93594 35600 93596
rect 35656 93594 35680 93596
rect 35736 93594 35760 93596
rect 35816 93594 35840 93596
rect 35896 93594 35902 93596
rect 35656 93542 35658 93594
rect 35838 93542 35840 93594
rect 35594 93540 35600 93542
rect 35656 93540 35680 93542
rect 35736 93540 35760 93542
rect 35816 93540 35840 93542
rect 35896 93540 35902 93542
rect 35594 93531 35902 93540
rect 4214 93052 4522 93061
rect 4214 93050 4220 93052
rect 4276 93050 4300 93052
rect 4356 93050 4380 93052
rect 4436 93050 4460 93052
rect 4516 93050 4522 93052
rect 4276 92998 4278 93050
rect 4458 92998 4460 93050
rect 4214 92996 4220 92998
rect 4276 92996 4300 92998
rect 4356 92996 4380 92998
rect 4436 92996 4460 92998
rect 4516 92996 4522 92998
rect 4214 92987 4522 92996
rect 34934 93052 35242 93061
rect 34934 93050 34940 93052
rect 34996 93050 35020 93052
rect 35076 93050 35100 93052
rect 35156 93050 35180 93052
rect 35236 93050 35242 93052
rect 34996 92998 34998 93050
rect 35178 92998 35180 93050
rect 34934 92996 34940 92998
rect 34996 92996 35020 92998
rect 35076 92996 35100 92998
rect 35156 92996 35180 92998
rect 35236 92996 35242 92998
rect 34934 92987 35242 92996
rect 4874 92508 5182 92517
rect 4874 92506 4880 92508
rect 4936 92506 4960 92508
rect 5016 92506 5040 92508
rect 5096 92506 5120 92508
rect 5176 92506 5182 92508
rect 4936 92454 4938 92506
rect 5118 92454 5120 92506
rect 4874 92452 4880 92454
rect 4936 92452 4960 92454
rect 5016 92452 5040 92454
rect 5096 92452 5120 92454
rect 5176 92452 5182 92454
rect 4874 92443 5182 92452
rect 35594 92508 35902 92517
rect 35594 92506 35600 92508
rect 35656 92506 35680 92508
rect 35736 92506 35760 92508
rect 35816 92506 35840 92508
rect 35896 92506 35902 92508
rect 35656 92454 35658 92506
rect 35838 92454 35840 92506
rect 35594 92452 35600 92454
rect 35656 92452 35680 92454
rect 35736 92452 35760 92454
rect 35816 92452 35840 92454
rect 35896 92452 35902 92454
rect 35594 92443 35902 92452
rect 4214 91964 4522 91973
rect 4214 91962 4220 91964
rect 4276 91962 4300 91964
rect 4356 91962 4380 91964
rect 4436 91962 4460 91964
rect 4516 91962 4522 91964
rect 4276 91910 4278 91962
rect 4458 91910 4460 91962
rect 4214 91908 4220 91910
rect 4276 91908 4300 91910
rect 4356 91908 4380 91910
rect 4436 91908 4460 91910
rect 4516 91908 4522 91910
rect 4214 91899 4522 91908
rect 34934 91964 35242 91973
rect 34934 91962 34940 91964
rect 34996 91962 35020 91964
rect 35076 91962 35100 91964
rect 35156 91962 35180 91964
rect 35236 91962 35242 91964
rect 34996 91910 34998 91962
rect 35178 91910 35180 91962
rect 34934 91908 34940 91910
rect 34996 91908 35020 91910
rect 35076 91908 35100 91910
rect 35156 91908 35180 91910
rect 35236 91908 35242 91910
rect 34934 91899 35242 91908
rect 4874 91420 5182 91429
rect 4874 91418 4880 91420
rect 4936 91418 4960 91420
rect 5016 91418 5040 91420
rect 5096 91418 5120 91420
rect 5176 91418 5182 91420
rect 4936 91366 4938 91418
rect 5118 91366 5120 91418
rect 4874 91364 4880 91366
rect 4936 91364 4960 91366
rect 5016 91364 5040 91366
rect 5096 91364 5120 91366
rect 5176 91364 5182 91366
rect 4874 91355 5182 91364
rect 35594 91420 35902 91429
rect 35594 91418 35600 91420
rect 35656 91418 35680 91420
rect 35736 91418 35760 91420
rect 35816 91418 35840 91420
rect 35896 91418 35902 91420
rect 35656 91366 35658 91418
rect 35838 91366 35840 91418
rect 35594 91364 35600 91366
rect 35656 91364 35680 91366
rect 35736 91364 35760 91366
rect 35816 91364 35840 91366
rect 35896 91364 35902 91366
rect 35594 91355 35902 91364
rect 4214 90876 4522 90885
rect 4214 90874 4220 90876
rect 4276 90874 4300 90876
rect 4356 90874 4380 90876
rect 4436 90874 4460 90876
rect 4516 90874 4522 90876
rect 4276 90822 4278 90874
rect 4458 90822 4460 90874
rect 4214 90820 4220 90822
rect 4276 90820 4300 90822
rect 4356 90820 4380 90822
rect 4436 90820 4460 90822
rect 4516 90820 4522 90822
rect 4214 90811 4522 90820
rect 34934 90876 35242 90885
rect 34934 90874 34940 90876
rect 34996 90874 35020 90876
rect 35076 90874 35100 90876
rect 35156 90874 35180 90876
rect 35236 90874 35242 90876
rect 34996 90822 34998 90874
rect 35178 90822 35180 90874
rect 34934 90820 34940 90822
rect 34996 90820 35020 90822
rect 35076 90820 35100 90822
rect 35156 90820 35180 90822
rect 35236 90820 35242 90822
rect 34934 90811 35242 90820
rect 4874 90332 5182 90341
rect 4874 90330 4880 90332
rect 4936 90330 4960 90332
rect 5016 90330 5040 90332
rect 5096 90330 5120 90332
rect 5176 90330 5182 90332
rect 4936 90278 4938 90330
rect 5118 90278 5120 90330
rect 4874 90276 4880 90278
rect 4936 90276 4960 90278
rect 5016 90276 5040 90278
rect 5096 90276 5120 90278
rect 5176 90276 5182 90278
rect 4874 90267 5182 90276
rect 35594 90332 35902 90341
rect 35594 90330 35600 90332
rect 35656 90330 35680 90332
rect 35736 90330 35760 90332
rect 35816 90330 35840 90332
rect 35896 90330 35902 90332
rect 35656 90278 35658 90330
rect 35838 90278 35840 90330
rect 35594 90276 35600 90278
rect 35656 90276 35680 90278
rect 35736 90276 35760 90278
rect 35816 90276 35840 90278
rect 35896 90276 35902 90278
rect 35594 90267 35902 90276
rect 4214 89788 4522 89797
rect 4214 89786 4220 89788
rect 4276 89786 4300 89788
rect 4356 89786 4380 89788
rect 4436 89786 4460 89788
rect 4516 89786 4522 89788
rect 4276 89734 4278 89786
rect 4458 89734 4460 89786
rect 4214 89732 4220 89734
rect 4276 89732 4300 89734
rect 4356 89732 4380 89734
rect 4436 89732 4460 89734
rect 4516 89732 4522 89734
rect 4214 89723 4522 89732
rect 34934 89788 35242 89797
rect 34934 89786 34940 89788
rect 34996 89786 35020 89788
rect 35076 89786 35100 89788
rect 35156 89786 35180 89788
rect 35236 89786 35242 89788
rect 34996 89734 34998 89786
rect 35178 89734 35180 89786
rect 34934 89732 34940 89734
rect 34996 89732 35020 89734
rect 35076 89732 35100 89734
rect 35156 89732 35180 89734
rect 35236 89732 35242 89734
rect 34934 89723 35242 89732
rect 4874 89244 5182 89253
rect 4874 89242 4880 89244
rect 4936 89242 4960 89244
rect 5016 89242 5040 89244
rect 5096 89242 5120 89244
rect 5176 89242 5182 89244
rect 4936 89190 4938 89242
rect 5118 89190 5120 89242
rect 4874 89188 4880 89190
rect 4936 89188 4960 89190
rect 5016 89188 5040 89190
rect 5096 89188 5120 89190
rect 5176 89188 5182 89190
rect 4874 89179 5182 89188
rect 35594 89244 35902 89253
rect 35594 89242 35600 89244
rect 35656 89242 35680 89244
rect 35736 89242 35760 89244
rect 35816 89242 35840 89244
rect 35896 89242 35902 89244
rect 35656 89190 35658 89242
rect 35838 89190 35840 89242
rect 35594 89188 35600 89190
rect 35656 89188 35680 89190
rect 35736 89188 35760 89190
rect 35816 89188 35840 89190
rect 35896 89188 35902 89190
rect 35594 89179 35902 89188
rect 4214 88700 4522 88709
rect 4214 88698 4220 88700
rect 4276 88698 4300 88700
rect 4356 88698 4380 88700
rect 4436 88698 4460 88700
rect 4516 88698 4522 88700
rect 4276 88646 4278 88698
rect 4458 88646 4460 88698
rect 4214 88644 4220 88646
rect 4276 88644 4300 88646
rect 4356 88644 4380 88646
rect 4436 88644 4460 88646
rect 4516 88644 4522 88646
rect 4214 88635 4522 88644
rect 34934 88700 35242 88709
rect 34934 88698 34940 88700
rect 34996 88698 35020 88700
rect 35076 88698 35100 88700
rect 35156 88698 35180 88700
rect 35236 88698 35242 88700
rect 34996 88646 34998 88698
rect 35178 88646 35180 88698
rect 34934 88644 34940 88646
rect 34996 88644 35020 88646
rect 35076 88644 35100 88646
rect 35156 88644 35180 88646
rect 35236 88644 35242 88646
rect 34934 88635 35242 88644
rect 4874 88156 5182 88165
rect 4874 88154 4880 88156
rect 4936 88154 4960 88156
rect 5016 88154 5040 88156
rect 5096 88154 5120 88156
rect 5176 88154 5182 88156
rect 4936 88102 4938 88154
rect 5118 88102 5120 88154
rect 4874 88100 4880 88102
rect 4936 88100 4960 88102
rect 5016 88100 5040 88102
rect 5096 88100 5120 88102
rect 5176 88100 5182 88102
rect 4874 88091 5182 88100
rect 35594 88156 35902 88165
rect 35594 88154 35600 88156
rect 35656 88154 35680 88156
rect 35736 88154 35760 88156
rect 35816 88154 35840 88156
rect 35896 88154 35902 88156
rect 35656 88102 35658 88154
rect 35838 88102 35840 88154
rect 35594 88100 35600 88102
rect 35656 88100 35680 88102
rect 35736 88100 35760 88102
rect 35816 88100 35840 88102
rect 35896 88100 35902 88102
rect 35594 88091 35902 88100
rect 4214 87612 4522 87621
rect 4214 87610 4220 87612
rect 4276 87610 4300 87612
rect 4356 87610 4380 87612
rect 4436 87610 4460 87612
rect 4516 87610 4522 87612
rect 4276 87558 4278 87610
rect 4458 87558 4460 87610
rect 4214 87556 4220 87558
rect 4276 87556 4300 87558
rect 4356 87556 4380 87558
rect 4436 87556 4460 87558
rect 4516 87556 4522 87558
rect 4214 87547 4522 87556
rect 34934 87612 35242 87621
rect 34934 87610 34940 87612
rect 34996 87610 35020 87612
rect 35076 87610 35100 87612
rect 35156 87610 35180 87612
rect 35236 87610 35242 87612
rect 34996 87558 34998 87610
rect 35178 87558 35180 87610
rect 34934 87556 34940 87558
rect 34996 87556 35020 87558
rect 35076 87556 35100 87558
rect 35156 87556 35180 87558
rect 35236 87556 35242 87558
rect 34934 87547 35242 87556
rect 4874 87068 5182 87077
rect 4874 87066 4880 87068
rect 4936 87066 4960 87068
rect 5016 87066 5040 87068
rect 5096 87066 5120 87068
rect 5176 87066 5182 87068
rect 4936 87014 4938 87066
rect 5118 87014 5120 87066
rect 4874 87012 4880 87014
rect 4936 87012 4960 87014
rect 5016 87012 5040 87014
rect 5096 87012 5120 87014
rect 5176 87012 5182 87014
rect 4874 87003 5182 87012
rect 35594 87068 35902 87077
rect 35594 87066 35600 87068
rect 35656 87066 35680 87068
rect 35736 87066 35760 87068
rect 35816 87066 35840 87068
rect 35896 87066 35902 87068
rect 35656 87014 35658 87066
rect 35838 87014 35840 87066
rect 35594 87012 35600 87014
rect 35656 87012 35680 87014
rect 35736 87012 35760 87014
rect 35816 87012 35840 87014
rect 35896 87012 35902 87014
rect 35594 87003 35902 87012
rect 4214 86524 4522 86533
rect 4214 86522 4220 86524
rect 4276 86522 4300 86524
rect 4356 86522 4380 86524
rect 4436 86522 4460 86524
rect 4516 86522 4522 86524
rect 4276 86470 4278 86522
rect 4458 86470 4460 86522
rect 4214 86468 4220 86470
rect 4276 86468 4300 86470
rect 4356 86468 4380 86470
rect 4436 86468 4460 86470
rect 4516 86468 4522 86470
rect 4214 86459 4522 86468
rect 34934 86524 35242 86533
rect 34934 86522 34940 86524
rect 34996 86522 35020 86524
rect 35076 86522 35100 86524
rect 35156 86522 35180 86524
rect 35236 86522 35242 86524
rect 34996 86470 34998 86522
rect 35178 86470 35180 86522
rect 34934 86468 34940 86470
rect 34996 86468 35020 86470
rect 35076 86468 35100 86470
rect 35156 86468 35180 86470
rect 35236 86468 35242 86470
rect 34934 86459 35242 86468
rect 4874 85980 5182 85989
rect 4874 85978 4880 85980
rect 4936 85978 4960 85980
rect 5016 85978 5040 85980
rect 5096 85978 5120 85980
rect 5176 85978 5182 85980
rect 4936 85926 4938 85978
rect 5118 85926 5120 85978
rect 4874 85924 4880 85926
rect 4936 85924 4960 85926
rect 5016 85924 5040 85926
rect 5096 85924 5120 85926
rect 5176 85924 5182 85926
rect 4874 85915 5182 85924
rect 35594 85980 35902 85989
rect 35594 85978 35600 85980
rect 35656 85978 35680 85980
rect 35736 85978 35760 85980
rect 35816 85978 35840 85980
rect 35896 85978 35902 85980
rect 35656 85926 35658 85978
rect 35838 85926 35840 85978
rect 35594 85924 35600 85926
rect 35656 85924 35680 85926
rect 35736 85924 35760 85926
rect 35816 85924 35840 85926
rect 35896 85924 35902 85926
rect 35594 85915 35902 85924
rect 4214 85436 4522 85445
rect 4214 85434 4220 85436
rect 4276 85434 4300 85436
rect 4356 85434 4380 85436
rect 4436 85434 4460 85436
rect 4516 85434 4522 85436
rect 4276 85382 4278 85434
rect 4458 85382 4460 85434
rect 4214 85380 4220 85382
rect 4276 85380 4300 85382
rect 4356 85380 4380 85382
rect 4436 85380 4460 85382
rect 4516 85380 4522 85382
rect 4214 85371 4522 85380
rect 34934 85436 35242 85445
rect 34934 85434 34940 85436
rect 34996 85434 35020 85436
rect 35076 85434 35100 85436
rect 35156 85434 35180 85436
rect 35236 85434 35242 85436
rect 34996 85382 34998 85434
rect 35178 85382 35180 85434
rect 34934 85380 34940 85382
rect 34996 85380 35020 85382
rect 35076 85380 35100 85382
rect 35156 85380 35180 85382
rect 35236 85380 35242 85382
rect 34934 85371 35242 85380
rect 4874 84892 5182 84901
rect 4874 84890 4880 84892
rect 4936 84890 4960 84892
rect 5016 84890 5040 84892
rect 5096 84890 5120 84892
rect 5176 84890 5182 84892
rect 4936 84838 4938 84890
rect 5118 84838 5120 84890
rect 4874 84836 4880 84838
rect 4936 84836 4960 84838
rect 5016 84836 5040 84838
rect 5096 84836 5120 84838
rect 5176 84836 5182 84838
rect 4874 84827 5182 84836
rect 35594 84892 35902 84901
rect 35594 84890 35600 84892
rect 35656 84890 35680 84892
rect 35736 84890 35760 84892
rect 35816 84890 35840 84892
rect 35896 84890 35902 84892
rect 35656 84838 35658 84890
rect 35838 84838 35840 84890
rect 35594 84836 35600 84838
rect 35656 84836 35680 84838
rect 35736 84836 35760 84838
rect 35816 84836 35840 84838
rect 35896 84836 35902 84838
rect 35594 84827 35902 84836
rect 4214 84348 4522 84357
rect 4214 84346 4220 84348
rect 4276 84346 4300 84348
rect 4356 84346 4380 84348
rect 4436 84346 4460 84348
rect 4516 84346 4522 84348
rect 4276 84294 4278 84346
rect 4458 84294 4460 84346
rect 4214 84292 4220 84294
rect 4276 84292 4300 84294
rect 4356 84292 4380 84294
rect 4436 84292 4460 84294
rect 4516 84292 4522 84294
rect 4214 84283 4522 84292
rect 34934 84348 35242 84357
rect 34934 84346 34940 84348
rect 34996 84346 35020 84348
rect 35076 84346 35100 84348
rect 35156 84346 35180 84348
rect 35236 84346 35242 84348
rect 34996 84294 34998 84346
rect 35178 84294 35180 84346
rect 34934 84292 34940 84294
rect 34996 84292 35020 84294
rect 35076 84292 35100 84294
rect 35156 84292 35180 84294
rect 35236 84292 35242 84294
rect 34934 84283 35242 84292
rect 4874 83804 5182 83813
rect 4874 83802 4880 83804
rect 4936 83802 4960 83804
rect 5016 83802 5040 83804
rect 5096 83802 5120 83804
rect 5176 83802 5182 83804
rect 4936 83750 4938 83802
rect 5118 83750 5120 83802
rect 4874 83748 4880 83750
rect 4936 83748 4960 83750
rect 5016 83748 5040 83750
rect 5096 83748 5120 83750
rect 5176 83748 5182 83750
rect 4874 83739 5182 83748
rect 35594 83804 35902 83813
rect 35594 83802 35600 83804
rect 35656 83802 35680 83804
rect 35736 83802 35760 83804
rect 35816 83802 35840 83804
rect 35896 83802 35902 83804
rect 35656 83750 35658 83802
rect 35838 83750 35840 83802
rect 35594 83748 35600 83750
rect 35656 83748 35680 83750
rect 35736 83748 35760 83750
rect 35816 83748 35840 83750
rect 35896 83748 35902 83750
rect 35594 83739 35902 83748
rect 4214 83260 4522 83269
rect 4214 83258 4220 83260
rect 4276 83258 4300 83260
rect 4356 83258 4380 83260
rect 4436 83258 4460 83260
rect 4516 83258 4522 83260
rect 4276 83206 4278 83258
rect 4458 83206 4460 83258
rect 4214 83204 4220 83206
rect 4276 83204 4300 83206
rect 4356 83204 4380 83206
rect 4436 83204 4460 83206
rect 4516 83204 4522 83206
rect 4214 83195 4522 83204
rect 34934 83260 35242 83269
rect 34934 83258 34940 83260
rect 34996 83258 35020 83260
rect 35076 83258 35100 83260
rect 35156 83258 35180 83260
rect 35236 83258 35242 83260
rect 34996 83206 34998 83258
rect 35178 83206 35180 83258
rect 34934 83204 34940 83206
rect 34996 83204 35020 83206
rect 35076 83204 35100 83206
rect 35156 83204 35180 83206
rect 35236 83204 35242 83206
rect 34934 83195 35242 83204
rect 4874 82716 5182 82725
rect 4874 82714 4880 82716
rect 4936 82714 4960 82716
rect 5016 82714 5040 82716
rect 5096 82714 5120 82716
rect 5176 82714 5182 82716
rect 4936 82662 4938 82714
rect 5118 82662 5120 82714
rect 4874 82660 4880 82662
rect 4936 82660 4960 82662
rect 5016 82660 5040 82662
rect 5096 82660 5120 82662
rect 5176 82660 5182 82662
rect 4874 82651 5182 82660
rect 35594 82716 35902 82725
rect 35594 82714 35600 82716
rect 35656 82714 35680 82716
rect 35736 82714 35760 82716
rect 35816 82714 35840 82716
rect 35896 82714 35902 82716
rect 35656 82662 35658 82714
rect 35838 82662 35840 82714
rect 35594 82660 35600 82662
rect 35656 82660 35680 82662
rect 35736 82660 35760 82662
rect 35816 82660 35840 82662
rect 35896 82660 35902 82662
rect 35594 82651 35902 82660
rect 4214 82172 4522 82181
rect 4214 82170 4220 82172
rect 4276 82170 4300 82172
rect 4356 82170 4380 82172
rect 4436 82170 4460 82172
rect 4516 82170 4522 82172
rect 4276 82118 4278 82170
rect 4458 82118 4460 82170
rect 4214 82116 4220 82118
rect 4276 82116 4300 82118
rect 4356 82116 4380 82118
rect 4436 82116 4460 82118
rect 4516 82116 4522 82118
rect 4214 82107 4522 82116
rect 34934 82172 35242 82181
rect 34934 82170 34940 82172
rect 34996 82170 35020 82172
rect 35076 82170 35100 82172
rect 35156 82170 35180 82172
rect 35236 82170 35242 82172
rect 34996 82118 34998 82170
rect 35178 82118 35180 82170
rect 34934 82116 34940 82118
rect 34996 82116 35020 82118
rect 35076 82116 35100 82118
rect 35156 82116 35180 82118
rect 35236 82116 35242 82118
rect 34934 82107 35242 82116
rect 4874 81628 5182 81637
rect 4874 81626 4880 81628
rect 4936 81626 4960 81628
rect 5016 81626 5040 81628
rect 5096 81626 5120 81628
rect 5176 81626 5182 81628
rect 4936 81574 4938 81626
rect 5118 81574 5120 81626
rect 4874 81572 4880 81574
rect 4936 81572 4960 81574
rect 5016 81572 5040 81574
rect 5096 81572 5120 81574
rect 5176 81572 5182 81574
rect 4874 81563 5182 81572
rect 35594 81628 35902 81637
rect 35594 81626 35600 81628
rect 35656 81626 35680 81628
rect 35736 81626 35760 81628
rect 35816 81626 35840 81628
rect 35896 81626 35902 81628
rect 35656 81574 35658 81626
rect 35838 81574 35840 81626
rect 35594 81572 35600 81574
rect 35656 81572 35680 81574
rect 35736 81572 35760 81574
rect 35816 81572 35840 81574
rect 35896 81572 35902 81574
rect 35594 81563 35902 81572
rect 4214 81084 4522 81093
rect 4214 81082 4220 81084
rect 4276 81082 4300 81084
rect 4356 81082 4380 81084
rect 4436 81082 4460 81084
rect 4516 81082 4522 81084
rect 4276 81030 4278 81082
rect 4458 81030 4460 81082
rect 4214 81028 4220 81030
rect 4276 81028 4300 81030
rect 4356 81028 4380 81030
rect 4436 81028 4460 81030
rect 4516 81028 4522 81030
rect 4214 81019 4522 81028
rect 34934 81084 35242 81093
rect 34934 81082 34940 81084
rect 34996 81082 35020 81084
rect 35076 81082 35100 81084
rect 35156 81082 35180 81084
rect 35236 81082 35242 81084
rect 34996 81030 34998 81082
rect 35178 81030 35180 81082
rect 34934 81028 34940 81030
rect 34996 81028 35020 81030
rect 35076 81028 35100 81030
rect 35156 81028 35180 81030
rect 35236 81028 35242 81030
rect 34934 81019 35242 81028
rect 4874 80540 5182 80549
rect 4874 80538 4880 80540
rect 4936 80538 4960 80540
rect 5016 80538 5040 80540
rect 5096 80538 5120 80540
rect 5176 80538 5182 80540
rect 4936 80486 4938 80538
rect 5118 80486 5120 80538
rect 4874 80484 4880 80486
rect 4936 80484 4960 80486
rect 5016 80484 5040 80486
rect 5096 80484 5120 80486
rect 5176 80484 5182 80486
rect 4874 80475 5182 80484
rect 35594 80540 35902 80549
rect 35594 80538 35600 80540
rect 35656 80538 35680 80540
rect 35736 80538 35760 80540
rect 35816 80538 35840 80540
rect 35896 80538 35902 80540
rect 35656 80486 35658 80538
rect 35838 80486 35840 80538
rect 35594 80484 35600 80486
rect 35656 80484 35680 80486
rect 35736 80484 35760 80486
rect 35816 80484 35840 80486
rect 35896 80484 35902 80486
rect 35594 80475 35902 80484
rect 4214 79996 4522 80005
rect 4214 79994 4220 79996
rect 4276 79994 4300 79996
rect 4356 79994 4380 79996
rect 4436 79994 4460 79996
rect 4516 79994 4522 79996
rect 4276 79942 4278 79994
rect 4458 79942 4460 79994
rect 4214 79940 4220 79942
rect 4276 79940 4300 79942
rect 4356 79940 4380 79942
rect 4436 79940 4460 79942
rect 4516 79940 4522 79942
rect 4214 79931 4522 79940
rect 34934 79996 35242 80005
rect 34934 79994 34940 79996
rect 34996 79994 35020 79996
rect 35076 79994 35100 79996
rect 35156 79994 35180 79996
rect 35236 79994 35242 79996
rect 34996 79942 34998 79994
rect 35178 79942 35180 79994
rect 34934 79940 34940 79942
rect 34996 79940 35020 79942
rect 35076 79940 35100 79942
rect 35156 79940 35180 79942
rect 35236 79940 35242 79942
rect 34934 79931 35242 79940
rect 4874 79452 5182 79461
rect 4874 79450 4880 79452
rect 4936 79450 4960 79452
rect 5016 79450 5040 79452
rect 5096 79450 5120 79452
rect 5176 79450 5182 79452
rect 4936 79398 4938 79450
rect 5118 79398 5120 79450
rect 4874 79396 4880 79398
rect 4936 79396 4960 79398
rect 5016 79396 5040 79398
rect 5096 79396 5120 79398
rect 5176 79396 5182 79398
rect 4874 79387 5182 79396
rect 35594 79452 35902 79461
rect 35594 79450 35600 79452
rect 35656 79450 35680 79452
rect 35736 79450 35760 79452
rect 35816 79450 35840 79452
rect 35896 79450 35902 79452
rect 35656 79398 35658 79450
rect 35838 79398 35840 79450
rect 35594 79396 35600 79398
rect 35656 79396 35680 79398
rect 35736 79396 35760 79398
rect 35816 79396 35840 79398
rect 35896 79396 35902 79398
rect 35594 79387 35902 79396
rect 4214 78908 4522 78917
rect 4214 78906 4220 78908
rect 4276 78906 4300 78908
rect 4356 78906 4380 78908
rect 4436 78906 4460 78908
rect 4516 78906 4522 78908
rect 4276 78854 4278 78906
rect 4458 78854 4460 78906
rect 4214 78852 4220 78854
rect 4276 78852 4300 78854
rect 4356 78852 4380 78854
rect 4436 78852 4460 78854
rect 4516 78852 4522 78854
rect 4214 78843 4522 78852
rect 34934 78908 35242 78917
rect 34934 78906 34940 78908
rect 34996 78906 35020 78908
rect 35076 78906 35100 78908
rect 35156 78906 35180 78908
rect 35236 78906 35242 78908
rect 34996 78854 34998 78906
rect 35178 78854 35180 78906
rect 34934 78852 34940 78854
rect 34996 78852 35020 78854
rect 35076 78852 35100 78854
rect 35156 78852 35180 78854
rect 35236 78852 35242 78854
rect 34934 78843 35242 78852
rect 4874 78364 5182 78373
rect 4874 78362 4880 78364
rect 4936 78362 4960 78364
rect 5016 78362 5040 78364
rect 5096 78362 5120 78364
rect 5176 78362 5182 78364
rect 4936 78310 4938 78362
rect 5118 78310 5120 78362
rect 4874 78308 4880 78310
rect 4936 78308 4960 78310
rect 5016 78308 5040 78310
rect 5096 78308 5120 78310
rect 5176 78308 5182 78310
rect 4874 78299 5182 78308
rect 35594 78364 35902 78373
rect 35594 78362 35600 78364
rect 35656 78362 35680 78364
rect 35736 78362 35760 78364
rect 35816 78362 35840 78364
rect 35896 78362 35902 78364
rect 35656 78310 35658 78362
rect 35838 78310 35840 78362
rect 35594 78308 35600 78310
rect 35656 78308 35680 78310
rect 35736 78308 35760 78310
rect 35816 78308 35840 78310
rect 35896 78308 35902 78310
rect 35594 78299 35902 78308
rect 4214 77820 4522 77829
rect 4214 77818 4220 77820
rect 4276 77818 4300 77820
rect 4356 77818 4380 77820
rect 4436 77818 4460 77820
rect 4516 77818 4522 77820
rect 4276 77766 4278 77818
rect 4458 77766 4460 77818
rect 4214 77764 4220 77766
rect 4276 77764 4300 77766
rect 4356 77764 4380 77766
rect 4436 77764 4460 77766
rect 4516 77764 4522 77766
rect 4214 77755 4522 77764
rect 34934 77820 35242 77829
rect 34934 77818 34940 77820
rect 34996 77818 35020 77820
rect 35076 77818 35100 77820
rect 35156 77818 35180 77820
rect 35236 77818 35242 77820
rect 34996 77766 34998 77818
rect 35178 77766 35180 77818
rect 34934 77764 34940 77766
rect 34996 77764 35020 77766
rect 35076 77764 35100 77766
rect 35156 77764 35180 77766
rect 35236 77764 35242 77766
rect 34934 77755 35242 77764
rect 43548 77722 43576 101390
rect 43536 77716 43588 77722
rect 43536 77658 43588 77664
rect 43628 77580 43680 77586
rect 43628 77522 43680 77528
rect 41788 77376 41840 77382
rect 41788 77318 41840 77324
rect 4874 77276 5182 77285
rect 4874 77274 4880 77276
rect 4936 77274 4960 77276
rect 5016 77274 5040 77276
rect 5096 77274 5120 77276
rect 5176 77274 5182 77276
rect 4936 77222 4938 77274
rect 5118 77222 5120 77274
rect 4874 77220 4880 77222
rect 4936 77220 4960 77222
rect 5016 77220 5040 77222
rect 5096 77220 5120 77222
rect 5176 77220 5182 77222
rect 4874 77211 5182 77220
rect 35594 77276 35902 77285
rect 35594 77274 35600 77276
rect 35656 77274 35680 77276
rect 35736 77274 35760 77276
rect 35816 77274 35840 77276
rect 35896 77274 35902 77276
rect 35656 77222 35658 77274
rect 35838 77222 35840 77274
rect 35594 77220 35600 77222
rect 35656 77220 35680 77222
rect 35736 77220 35760 77222
rect 35816 77220 35840 77222
rect 35896 77220 35902 77222
rect 35594 77211 35902 77220
rect 41800 76838 41828 77318
rect 43640 77042 43668 77522
rect 45388 77178 45416 101390
rect 47504 77722 47532 101390
rect 49712 77722 49740 101390
rect 47492 77716 47544 77722
rect 47492 77658 47544 77664
rect 49700 77716 49752 77722
rect 49700 77658 49752 77664
rect 49424 77580 49476 77586
rect 49424 77522 49476 77528
rect 45652 77444 45704 77450
rect 45652 77386 45704 77392
rect 45744 77444 45796 77450
rect 45744 77386 45796 77392
rect 47952 77444 48004 77450
rect 47952 77386 48004 77392
rect 45376 77172 45428 77178
rect 45376 77114 45428 77120
rect 43628 77036 43680 77042
rect 43628 76978 43680 76984
rect 43628 76900 43680 76906
rect 43628 76842 43680 76848
rect 41788 76832 41840 76838
rect 41788 76774 41840 76780
rect 4214 76732 4522 76741
rect 4214 76730 4220 76732
rect 4276 76730 4300 76732
rect 4356 76730 4380 76732
rect 4436 76730 4460 76732
rect 4516 76730 4522 76732
rect 4276 76678 4278 76730
rect 4458 76678 4460 76730
rect 4214 76676 4220 76678
rect 4276 76676 4300 76678
rect 4356 76676 4380 76678
rect 4436 76676 4460 76678
rect 4516 76676 4522 76678
rect 4214 76667 4522 76676
rect 34934 76732 35242 76741
rect 34934 76730 34940 76732
rect 34996 76730 35020 76732
rect 35076 76730 35100 76732
rect 35156 76730 35180 76732
rect 35236 76730 35242 76732
rect 34996 76678 34998 76730
rect 35178 76678 35180 76730
rect 34934 76676 34940 76678
rect 34996 76676 35020 76678
rect 35076 76676 35100 76678
rect 35156 76676 35180 76678
rect 35236 76676 35242 76678
rect 34934 76667 35242 76676
rect 4874 76188 5182 76197
rect 4874 76186 4880 76188
rect 4936 76186 4960 76188
rect 5016 76186 5040 76188
rect 5096 76186 5120 76188
rect 5176 76186 5182 76188
rect 4936 76134 4938 76186
rect 5118 76134 5120 76186
rect 4874 76132 4880 76134
rect 4936 76132 4960 76134
rect 5016 76132 5040 76134
rect 5096 76132 5120 76134
rect 5176 76132 5182 76134
rect 4874 76123 5182 76132
rect 35594 76188 35902 76197
rect 35594 76186 35600 76188
rect 35656 76186 35680 76188
rect 35736 76186 35760 76188
rect 35816 76186 35840 76188
rect 35896 76186 35902 76188
rect 35656 76134 35658 76186
rect 35838 76134 35840 76186
rect 35594 76132 35600 76134
rect 35656 76132 35680 76134
rect 35736 76132 35760 76134
rect 35816 76132 35840 76134
rect 35896 76132 35902 76134
rect 35594 76123 35902 76132
rect 4214 75644 4522 75653
rect 4214 75642 4220 75644
rect 4276 75642 4300 75644
rect 4356 75642 4380 75644
rect 4436 75642 4460 75644
rect 4516 75642 4522 75644
rect 4276 75590 4278 75642
rect 4458 75590 4460 75642
rect 4214 75588 4220 75590
rect 4276 75588 4300 75590
rect 4356 75588 4380 75590
rect 4436 75588 4460 75590
rect 4516 75588 4522 75590
rect 4214 75579 4522 75588
rect 34934 75644 35242 75653
rect 34934 75642 34940 75644
rect 34996 75642 35020 75644
rect 35076 75642 35100 75644
rect 35156 75642 35180 75644
rect 35236 75642 35242 75644
rect 34996 75590 34998 75642
rect 35178 75590 35180 75642
rect 34934 75588 34940 75590
rect 34996 75588 35020 75590
rect 35076 75588 35100 75590
rect 35156 75588 35180 75590
rect 35236 75588 35242 75590
rect 34934 75579 35242 75588
rect 4874 75100 5182 75109
rect 4874 75098 4880 75100
rect 4936 75098 4960 75100
rect 5016 75098 5040 75100
rect 5096 75098 5120 75100
rect 5176 75098 5182 75100
rect 4936 75046 4938 75098
rect 5118 75046 5120 75098
rect 4874 75044 4880 75046
rect 4936 75044 4960 75046
rect 5016 75044 5040 75046
rect 5096 75044 5120 75046
rect 5176 75044 5182 75046
rect 4874 75035 5182 75044
rect 35594 75100 35902 75109
rect 35594 75098 35600 75100
rect 35656 75098 35680 75100
rect 35736 75098 35760 75100
rect 35816 75098 35840 75100
rect 35896 75098 35902 75100
rect 35656 75046 35658 75098
rect 35838 75046 35840 75098
rect 35594 75044 35600 75046
rect 35656 75044 35680 75046
rect 35736 75044 35760 75046
rect 35816 75044 35840 75046
rect 35896 75044 35902 75046
rect 35594 75035 35902 75044
rect 4214 74556 4522 74565
rect 4214 74554 4220 74556
rect 4276 74554 4300 74556
rect 4356 74554 4380 74556
rect 4436 74554 4460 74556
rect 4516 74554 4522 74556
rect 4276 74502 4278 74554
rect 4458 74502 4460 74554
rect 4214 74500 4220 74502
rect 4276 74500 4300 74502
rect 4356 74500 4380 74502
rect 4436 74500 4460 74502
rect 4516 74500 4522 74502
rect 4214 74491 4522 74500
rect 34934 74556 35242 74565
rect 34934 74554 34940 74556
rect 34996 74554 35020 74556
rect 35076 74554 35100 74556
rect 35156 74554 35180 74556
rect 35236 74554 35242 74556
rect 34996 74502 34998 74554
rect 35178 74502 35180 74554
rect 34934 74500 34940 74502
rect 34996 74500 35020 74502
rect 35076 74500 35100 74502
rect 35156 74500 35180 74502
rect 35236 74500 35242 74502
rect 34934 74491 35242 74500
rect 4874 74012 5182 74021
rect 4874 74010 4880 74012
rect 4936 74010 4960 74012
rect 5016 74010 5040 74012
rect 5096 74010 5120 74012
rect 5176 74010 5182 74012
rect 4936 73958 4938 74010
rect 5118 73958 5120 74010
rect 4874 73956 4880 73958
rect 4936 73956 4960 73958
rect 5016 73956 5040 73958
rect 5096 73956 5120 73958
rect 5176 73956 5182 73958
rect 4874 73947 5182 73956
rect 35594 74012 35902 74021
rect 35594 74010 35600 74012
rect 35656 74010 35680 74012
rect 35736 74010 35760 74012
rect 35816 74010 35840 74012
rect 35896 74010 35902 74012
rect 35656 73958 35658 74010
rect 35838 73958 35840 74010
rect 35594 73956 35600 73958
rect 35656 73956 35680 73958
rect 35736 73956 35760 73958
rect 35816 73956 35840 73958
rect 35896 73956 35902 73958
rect 35594 73947 35902 73956
rect 4214 73468 4522 73477
rect 4214 73466 4220 73468
rect 4276 73466 4300 73468
rect 4356 73466 4380 73468
rect 4436 73466 4460 73468
rect 4516 73466 4522 73468
rect 4276 73414 4278 73466
rect 4458 73414 4460 73466
rect 4214 73412 4220 73414
rect 4276 73412 4300 73414
rect 4356 73412 4380 73414
rect 4436 73412 4460 73414
rect 4516 73412 4522 73414
rect 4214 73403 4522 73412
rect 34934 73468 35242 73477
rect 34934 73466 34940 73468
rect 34996 73466 35020 73468
rect 35076 73466 35100 73468
rect 35156 73466 35180 73468
rect 35236 73466 35242 73468
rect 34996 73414 34998 73466
rect 35178 73414 35180 73466
rect 34934 73412 34940 73414
rect 34996 73412 35020 73414
rect 35076 73412 35100 73414
rect 35156 73412 35180 73414
rect 35236 73412 35242 73414
rect 34934 73403 35242 73412
rect 4874 72924 5182 72933
rect 4874 72922 4880 72924
rect 4936 72922 4960 72924
rect 5016 72922 5040 72924
rect 5096 72922 5120 72924
rect 5176 72922 5182 72924
rect 4936 72870 4938 72922
rect 5118 72870 5120 72922
rect 4874 72868 4880 72870
rect 4936 72868 4960 72870
rect 5016 72868 5040 72870
rect 5096 72868 5120 72870
rect 5176 72868 5182 72870
rect 4874 72859 5182 72868
rect 35594 72924 35902 72933
rect 35594 72922 35600 72924
rect 35656 72922 35680 72924
rect 35736 72922 35760 72924
rect 35816 72922 35840 72924
rect 35896 72922 35902 72924
rect 35656 72870 35658 72922
rect 35838 72870 35840 72922
rect 35594 72868 35600 72870
rect 35656 72868 35680 72870
rect 35736 72868 35760 72870
rect 35816 72868 35840 72870
rect 35896 72868 35902 72870
rect 35594 72859 35902 72868
rect 4214 72380 4522 72389
rect 4214 72378 4220 72380
rect 4276 72378 4300 72380
rect 4356 72378 4380 72380
rect 4436 72378 4460 72380
rect 4516 72378 4522 72380
rect 4276 72326 4278 72378
rect 4458 72326 4460 72378
rect 4214 72324 4220 72326
rect 4276 72324 4300 72326
rect 4356 72324 4380 72326
rect 4436 72324 4460 72326
rect 4516 72324 4522 72326
rect 4214 72315 4522 72324
rect 34934 72380 35242 72389
rect 34934 72378 34940 72380
rect 34996 72378 35020 72380
rect 35076 72378 35100 72380
rect 35156 72378 35180 72380
rect 35236 72378 35242 72380
rect 34996 72326 34998 72378
rect 35178 72326 35180 72378
rect 34934 72324 34940 72326
rect 34996 72324 35020 72326
rect 35076 72324 35100 72326
rect 35156 72324 35180 72326
rect 35236 72324 35242 72326
rect 34934 72315 35242 72324
rect 4874 71836 5182 71845
rect 4874 71834 4880 71836
rect 4936 71834 4960 71836
rect 5016 71834 5040 71836
rect 5096 71834 5120 71836
rect 5176 71834 5182 71836
rect 4936 71782 4938 71834
rect 5118 71782 5120 71834
rect 4874 71780 4880 71782
rect 4936 71780 4960 71782
rect 5016 71780 5040 71782
rect 5096 71780 5120 71782
rect 5176 71780 5182 71782
rect 4874 71771 5182 71780
rect 35594 71836 35902 71845
rect 35594 71834 35600 71836
rect 35656 71834 35680 71836
rect 35736 71834 35760 71836
rect 35816 71834 35840 71836
rect 35896 71834 35902 71836
rect 35656 71782 35658 71834
rect 35838 71782 35840 71834
rect 35594 71780 35600 71782
rect 35656 71780 35680 71782
rect 35736 71780 35760 71782
rect 35816 71780 35840 71782
rect 35896 71780 35902 71782
rect 35594 71771 35902 71780
rect 4214 71292 4522 71301
rect 4214 71290 4220 71292
rect 4276 71290 4300 71292
rect 4356 71290 4380 71292
rect 4436 71290 4460 71292
rect 4516 71290 4522 71292
rect 4276 71238 4278 71290
rect 4458 71238 4460 71290
rect 4214 71236 4220 71238
rect 4276 71236 4300 71238
rect 4356 71236 4380 71238
rect 4436 71236 4460 71238
rect 4516 71236 4522 71238
rect 4214 71227 4522 71236
rect 34934 71292 35242 71301
rect 34934 71290 34940 71292
rect 34996 71290 35020 71292
rect 35076 71290 35100 71292
rect 35156 71290 35180 71292
rect 35236 71290 35242 71292
rect 34996 71238 34998 71290
rect 35178 71238 35180 71290
rect 34934 71236 34940 71238
rect 34996 71236 35020 71238
rect 35076 71236 35100 71238
rect 35156 71236 35180 71238
rect 35236 71236 35242 71238
rect 34934 71227 35242 71236
rect 4874 70748 5182 70757
rect 4874 70746 4880 70748
rect 4936 70746 4960 70748
rect 5016 70746 5040 70748
rect 5096 70746 5120 70748
rect 5176 70746 5182 70748
rect 4936 70694 4938 70746
rect 5118 70694 5120 70746
rect 4874 70692 4880 70694
rect 4936 70692 4960 70694
rect 5016 70692 5040 70694
rect 5096 70692 5120 70694
rect 5176 70692 5182 70694
rect 4874 70683 5182 70692
rect 35594 70748 35902 70757
rect 35594 70746 35600 70748
rect 35656 70746 35680 70748
rect 35736 70746 35760 70748
rect 35816 70746 35840 70748
rect 35896 70746 35902 70748
rect 35656 70694 35658 70746
rect 35838 70694 35840 70746
rect 35594 70692 35600 70694
rect 35656 70692 35680 70694
rect 35736 70692 35760 70694
rect 35816 70692 35840 70694
rect 35896 70692 35902 70694
rect 35594 70683 35902 70692
rect 4214 70204 4522 70213
rect 4214 70202 4220 70204
rect 4276 70202 4300 70204
rect 4356 70202 4380 70204
rect 4436 70202 4460 70204
rect 4516 70202 4522 70204
rect 4276 70150 4278 70202
rect 4458 70150 4460 70202
rect 4214 70148 4220 70150
rect 4276 70148 4300 70150
rect 4356 70148 4380 70150
rect 4436 70148 4460 70150
rect 4516 70148 4522 70150
rect 4214 70139 4522 70148
rect 34934 70204 35242 70213
rect 34934 70202 34940 70204
rect 34996 70202 35020 70204
rect 35076 70202 35100 70204
rect 35156 70202 35180 70204
rect 35236 70202 35242 70204
rect 34996 70150 34998 70202
rect 35178 70150 35180 70202
rect 34934 70148 34940 70150
rect 34996 70148 35020 70150
rect 35076 70148 35100 70150
rect 35156 70148 35180 70150
rect 35236 70148 35242 70150
rect 34934 70139 35242 70148
rect 4874 69660 5182 69669
rect 4874 69658 4880 69660
rect 4936 69658 4960 69660
rect 5016 69658 5040 69660
rect 5096 69658 5120 69660
rect 5176 69658 5182 69660
rect 4936 69606 4938 69658
rect 5118 69606 5120 69658
rect 4874 69604 4880 69606
rect 4936 69604 4960 69606
rect 5016 69604 5040 69606
rect 5096 69604 5120 69606
rect 5176 69604 5182 69606
rect 4874 69595 5182 69604
rect 35594 69660 35902 69669
rect 35594 69658 35600 69660
rect 35656 69658 35680 69660
rect 35736 69658 35760 69660
rect 35816 69658 35840 69660
rect 35896 69658 35902 69660
rect 35656 69606 35658 69658
rect 35838 69606 35840 69658
rect 35594 69604 35600 69606
rect 35656 69604 35680 69606
rect 35736 69604 35760 69606
rect 35816 69604 35840 69606
rect 35896 69604 35902 69606
rect 35594 69595 35902 69604
rect 4214 69116 4522 69125
rect 4214 69114 4220 69116
rect 4276 69114 4300 69116
rect 4356 69114 4380 69116
rect 4436 69114 4460 69116
rect 4516 69114 4522 69116
rect 4276 69062 4278 69114
rect 4458 69062 4460 69114
rect 4214 69060 4220 69062
rect 4276 69060 4300 69062
rect 4356 69060 4380 69062
rect 4436 69060 4460 69062
rect 4516 69060 4522 69062
rect 4214 69051 4522 69060
rect 34934 69116 35242 69125
rect 34934 69114 34940 69116
rect 34996 69114 35020 69116
rect 35076 69114 35100 69116
rect 35156 69114 35180 69116
rect 35236 69114 35242 69116
rect 34996 69062 34998 69114
rect 35178 69062 35180 69114
rect 34934 69060 34940 69062
rect 34996 69060 35020 69062
rect 35076 69060 35100 69062
rect 35156 69060 35180 69062
rect 35236 69060 35242 69062
rect 34934 69051 35242 69060
rect 4874 68572 5182 68581
rect 4874 68570 4880 68572
rect 4936 68570 4960 68572
rect 5016 68570 5040 68572
rect 5096 68570 5120 68572
rect 5176 68570 5182 68572
rect 4936 68518 4938 68570
rect 5118 68518 5120 68570
rect 4874 68516 4880 68518
rect 4936 68516 4960 68518
rect 5016 68516 5040 68518
rect 5096 68516 5120 68518
rect 5176 68516 5182 68518
rect 4874 68507 5182 68516
rect 35594 68572 35902 68581
rect 35594 68570 35600 68572
rect 35656 68570 35680 68572
rect 35736 68570 35760 68572
rect 35816 68570 35840 68572
rect 35896 68570 35902 68572
rect 35656 68518 35658 68570
rect 35838 68518 35840 68570
rect 35594 68516 35600 68518
rect 35656 68516 35680 68518
rect 35736 68516 35760 68518
rect 35816 68516 35840 68518
rect 35896 68516 35902 68518
rect 35594 68507 35902 68516
rect 4214 68028 4522 68037
rect 4214 68026 4220 68028
rect 4276 68026 4300 68028
rect 4356 68026 4380 68028
rect 4436 68026 4460 68028
rect 4516 68026 4522 68028
rect 4276 67974 4278 68026
rect 4458 67974 4460 68026
rect 4214 67972 4220 67974
rect 4276 67972 4300 67974
rect 4356 67972 4380 67974
rect 4436 67972 4460 67974
rect 4516 67972 4522 67974
rect 4214 67963 4522 67972
rect 34934 68028 35242 68037
rect 34934 68026 34940 68028
rect 34996 68026 35020 68028
rect 35076 68026 35100 68028
rect 35156 68026 35180 68028
rect 35236 68026 35242 68028
rect 34996 67974 34998 68026
rect 35178 67974 35180 68026
rect 34934 67972 34940 67974
rect 34996 67972 35020 67974
rect 35076 67972 35100 67974
rect 35156 67972 35180 67974
rect 35236 67972 35242 67974
rect 34934 67963 35242 67972
rect 4874 67484 5182 67493
rect 4874 67482 4880 67484
rect 4936 67482 4960 67484
rect 5016 67482 5040 67484
rect 5096 67482 5120 67484
rect 5176 67482 5182 67484
rect 4936 67430 4938 67482
rect 5118 67430 5120 67482
rect 4874 67428 4880 67430
rect 4936 67428 4960 67430
rect 5016 67428 5040 67430
rect 5096 67428 5120 67430
rect 5176 67428 5182 67430
rect 4874 67419 5182 67428
rect 35594 67484 35902 67493
rect 35594 67482 35600 67484
rect 35656 67482 35680 67484
rect 35736 67482 35760 67484
rect 35816 67482 35840 67484
rect 35896 67482 35902 67484
rect 35656 67430 35658 67482
rect 35838 67430 35840 67482
rect 35594 67428 35600 67430
rect 35656 67428 35680 67430
rect 35736 67428 35760 67430
rect 35816 67428 35840 67430
rect 35896 67428 35902 67430
rect 35594 67419 35902 67428
rect 4214 66940 4522 66949
rect 4214 66938 4220 66940
rect 4276 66938 4300 66940
rect 4356 66938 4380 66940
rect 4436 66938 4460 66940
rect 4516 66938 4522 66940
rect 4276 66886 4278 66938
rect 4458 66886 4460 66938
rect 4214 66884 4220 66886
rect 4276 66884 4300 66886
rect 4356 66884 4380 66886
rect 4436 66884 4460 66886
rect 4516 66884 4522 66886
rect 4214 66875 4522 66884
rect 34934 66940 35242 66949
rect 34934 66938 34940 66940
rect 34996 66938 35020 66940
rect 35076 66938 35100 66940
rect 35156 66938 35180 66940
rect 35236 66938 35242 66940
rect 34996 66886 34998 66938
rect 35178 66886 35180 66938
rect 34934 66884 34940 66886
rect 34996 66884 35020 66886
rect 35076 66884 35100 66886
rect 35156 66884 35180 66886
rect 35236 66884 35242 66886
rect 34934 66875 35242 66884
rect 4874 66396 5182 66405
rect 4874 66394 4880 66396
rect 4936 66394 4960 66396
rect 5016 66394 5040 66396
rect 5096 66394 5120 66396
rect 5176 66394 5182 66396
rect 4936 66342 4938 66394
rect 5118 66342 5120 66394
rect 4874 66340 4880 66342
rect 4936 66340 4960 66342
rect 5016 66340 5040 66342
rect 5096 66340 5120 66342
rect 5176 66340 5182 66342
rect 4874 66331 5182 66340
rect 35594 66396 35902 66405
rect 35594 66394 35600 66396
rect 35656 66394 35680 66396
rect 35736 66394 35760 66396
rect 35816 66394 35840 66396
rect 35896 66394 35902 66396
rect 35656 66342 35658 66394
rect 35838 66342 35840 66394
rect 35594 66340 35600 66342
rect 35656 66340 35680 66342
rect 35736 66340 35760 66342
rect 35816 66340 35840 66342
rect 35896 66340 35902 66342
rect 35594 66331 35902 66340
rect 4214 65852 4522 65861
rect 4214 65850 4220 65852
rect 4276 65850 4300 65852
rect 4356 65850 4380 65852
rect 4436 65850 4460 65852
rect 4516 65850 4522 65852
rect 4276 65798 4278 65850
rect 4458 65798 4460 65850
rect 4214 65796 4220 65798
rect 4276 65796 4300 65798
rect 4356 65796 4380 65798
rect 4436 65796 4460 65798
rect 4516 65796 4522 65798
rect 4214 65787 4522 65796
rect 34934 65852 35242 65861
rect 34934 65850 34940 65852
rect 34996 65850 35020 65852
rect 35076 65850 35100 65852
rect 35156 65850 35180 65852
rect 35236 65850 35242 65852
rect 34996 65798 34998 65850
rect 35178 65798 35180 65850
rect 34934 65796 34940 65798
rect 34996 65796 35020 65798
rect 35076 65796 35100 65798
rect 35156 65796 35180 65798
rect 35236 65796 35242 65798
rect 34934 65787 35242 65796
rect 4874 65308 5182 65317
rect 4874 65306 4880 65308
rect 4936 65306 4960 65308
rect 5016 65306 5040 65308
rect 5096 65306 5120 65308
rect 5176 65306 5182 65308
rect 4936 65254 4938 65306
rect 5118 65254 5120 65306
rect 4874 65252 4880 65254
rect 4936 65252 4960 65254
rect 5016 65252 5040 65254
rect 5096 65252 5120 65254
rect 5176 65252 5182 65254
rect 4874 65243 5182 65252
rect 35594 65308 35902 65317
rect 35594 65306 35600 65308
rect 35656 65306 35680 65308
rect 35736 65306 35760 65308
rect 35816 65306 35840 65308
rect 35896 65306 35902 65308
rect 35656 65254 35658 65306
rect 35838 65254 35840 65306
rect 35594 65252 35600 65254
rect 35656 65252 35680 65254
rect 35736 65252 35760 65254
rect 35816 65252 35840 65254
rect 35896 65252 35902 65254
rect 35594 65243 35902 65252
rect 4214 64764 4522 64773
rect 4214 64762 4220 64764
rect 4276 64762 4300 64764
rect 4356 64762 4380 64764
rect 4436 64762 4460 64764
rect 4516 64762 4522 64764
rect 4276 64710 4278 64762
rect 4458 64710 4460 64762
rect 4214 64708 4220 64710
rect 4276 64708 4300 64710
rect 4356 64708 4380 64710
rect 4436 64708 4460 64710
rect 4516 64708 4522 64710
rect 4214 64699 4522 64708
rect 34934 64764 35242 64773
rect 34934 64762 34940 64764
rect 34996 64762 35020 64764
rect 35076 64762 35100 64764
rect 35156 64762 35180 64764
rect 35236 64762 35242 64764
rect 34996 64710 34998 64762
rect 35178 64710 35180 64762
rect 34934 64708 34940 64710
rect 34996 64708 35020 64710
rect 35076 64708 35100 64710
rect 35156 64708 35180 64710
rect 35236 64708 35242 64710
rect 34934 64699 35242 64708
rect 4874 64220 5182 64229
rect 4874 64218 4880 64220
rect 4936 64218 4960 64220
rect 5016 64218 5040 64220
rect 5096 64218 5120 64220
rect 5176 64218 5182 64220
rect 4936 64166 4938 64218
rect 5118 64166 5120 64218
rect 4874 64164 4880 64166
rect 4936 64164 4960 64166
rect 5016 64164 5040 64166
rect 5096 64164 5120 64166
rect 5176 64164 5182 64166
rect 4874 64155 5182 64164
rect 35594 64220 35902 64229
rect 35594 64218 35600 64220
rect 35656 64218 35680 64220
rect 35736 64218 35760 64220
rect 35816 64218 35840 64220
rect 35896 64218 35902 64220
rect 35656 64166 35658 64218
rect 35838 64166 35840 64218
rect 35594 64164 35600 64166
rect 35656 64164 35680 64166
rect 35736 64164 35760 64166
rect 35816 64164 35840 64166
rect 35896 64164 35902 64166
rect 35594 64155 35902 64164
rect 4214 63676 4522 63685
rect 4214 63674 4220 63676
rect 4276 63674 4300 63676
rect 4356 63674 4380 63676
rect 4436 63674 4460 63676
rect 4516 63674 4522 63676
rect 4276 63622 4278 63674
rect 4458 63622 4460 63674
rect 4214 63620 4220 63622
rect 4276 63620 4300 63622
rect 4356 63620 4380 63622
rect 4436 63620 4460 63622
rect 4516 63620 4522 63622
rect 4214 63611 4522 63620
rect 34934 63676 35242 63685
rect 34934 63674 34940 63676
rect 34996 63674 35020 63676
rect 35076 63674 35100 63676
rect 35156 63674 35180 63676
rect 35236 63674 35242 63676
rect 34996 63622 34998 63674
rect 35178 63622 35180 63674
rect 34934 63620 34940 63622
rect 34996 63620 35020 63622
rect 35076 63620 35100 63622
rect 35156 63620 35180 63622
rect 35236 63620 35242 63622
rect 34934 63611 35242 63620
rect 4874 63132 5182 63141
rect 4874 63130 4880 63132
rect 4936 63130 4960 63132
rect 5016 63130 5040 63132
rect 5096 63130 5120 63132
rect 5176 63130 5182 63132
rect 4936 63078 4938 63130
rect 5118 63078 5120 63130
rect 4874 63076 4880 63078
rect 4936 63076 4960 63078
rect 5016 63076 5040 63078
rect 5096 63076 5120 63078
rect 5176 63076 5182 63078
rect 4874 63067 5182 63076
rect 35594 63132 35902 63141
rect 35594 63130 35600 63132
rect 35656 63130 35680 63132
rect 35736 63130 35760 63132
rect 35816 63130 35840 63132
rect 35896 63130 35902 63132
rect 35656 63078 35658 63130
rect 35838 63078 35840 63130
rect 35594 63076 35600 63078
rect 35656 63076 35680 63078
rect 35736 63076 35760 63078
rect 35816 63076 35840 63078
rect 35896 63076 35902 63078
rect 35594 63067 35902 63076
rect 41800 62801 41828 76774
rect 43640 76294 43668 76842
rect 43628 76288 43680 76294
rect 43626 76256 43628 76265
rect 43680 76256 43682 76265
rect 43626 76191 43682 76200
rect 45664 75002 45692 77386
rect 45756 76838 45784 77386
rect 47964 76838 47992 77386
rect 48228 77104 48280 77110
rect 48228 77046 48280 77052
rect 45744 76832 45796 76838
rect 45744 76774 45796 76780
rect 47952 76832 48004 76838
rect 47952 76774 48004 76780
rect 45652 74996 45704 75002
rect 45652 74938 45704 74944
rect 45756 74633 45784 76774
rect 47964 75993 47992 76774
rect 47950 75984 48006 75993
rect 47950 75919 48006 75928
rect 48240 75002 48268 77046
rect 49436 77042 49464 77522
rect 51080 77444 51132 77450
rect 51080 77386 51132 77392
rect 49976 77376 50028 77382
rect 49976 77318 50028 77324
rect 49608 77104 49660 77110
rect 49606 77072 49608 77081
rect 49660 77072 49662 77081
rect 49424 77036 49476 77042
rect 49606 77007 49662 77016
rect 49424 76978 49476 76984
rect 48228 74996 48280 75002
rect 48228 74938 48280 74944
rect 46664 74860 46716 74866
rect 46664 74802 46716 74808
rect 45742 74624 45798 74633
rect 45742 74559 45798 74568
rect 41786 62792 41842 62801
rect 41786 62727 41842 62736
rect 4214 62588 4522 62597
rect 4214 62586 4220 62588
rect 4276 62586 4300 62588
rect 4356 62586 4380 62588
rect 4436 62586 4460 62588
rect 4516 62586 4522 62588
rect 4276 62534 4278 62586
rect 4458 62534 4460 62586
rect 4214 62532 4220 62534
rect 4276 62532 4300 62534
rect 4356 62532 4380 62534
rect 4436 62532 4460 62534
rect 4516 62532 4522 62534
rect 4214 62523 4522 62532
rect 34934 62588 35242 62597
rect 34934 62586 34940 62588
rect 34996 62586 35020 62588
rect 35076 62586 35100 62588
rect 35156 62586 35180 62588
rect 35236 62586 35242 62588
rect 34996 62534 34998 62586
rect 35178 62534 35180 62586
rect 34934 62532 34940 62534
rect 34996 62532 35020 62534
rect 35076 62532 35100 62534
rect 35156 62532 35180 62534
rect 35236 62532 35242 62534
rect 34934 62523 35242 62532
rect 1492 62144 1544 62150
rect 1492 62086 1544 62092
rect 1860 62144 1912 62150
rect 1860 62086 1912 62092
rect 1504 61985 1532 62086
rect 1490 61976 1546 61985
rect 1490 61911 1546 61920
rect 848 61600 900 61606
rect 848 61542 900 61548
rect 860 61441 888 61542
rect 846 61432 902 61441
rect 846 61367 902 61376
rect 1872 60518 1900 62086
rect 4874 62044 5182 62053
rect 4874 62042 4880 62044
rect 4936 62042 4960 62044
rect 5016 62042 5040 62044
rect 5096 62042 5120 62044
rect 5176 62042 5182 62044
rect 4936 61990 4938 62042
rect 5118 61990 5120 62042
rect 4874 61988 4880 61990
rect 4936 61988 4960 61990
rect 5016 61988 5040 61990
rect 5096 61988 5120 61990
rect 5176 61988 5182 61990
rect 4874 61979 5182 61988
rect 35594 62044 35902 62053
rect 35594 62042 35600 62044
rect 35656 62042 35680 62044
rect 35736 62042 35760 62044
rect 35816 62042 35840 62044
rect 35896 62042 35902 62044
rect 35656 61990 35658 62042
rect 35838 61990 35840 62042
rect 35594 61988 35600 61990
rect 35656 61988 35680 61990
rect 35736 61988 35760 61990
rect 35816 61988 35840 61990
rect 35896 61988 35902 61990
rect 35594 61979 35902 61988
rect 21088 61804 21140 61810
rect 21088 61746 21140 61752
rect 4214 61500 4522 61509
rect 4214 61498 4220 61500
rect 4276 61498 4300 61500
rect 4356 61498 4380 61500
rect 4436 61498 4460 61500
rect 4516 61498 4522 61500
rect 4276 61446 4278 61498
rect 4458 61446 4460 61498
rect 4214 61444 4220 61446
rect 4276 61444 4300 61446
rect 4356 61444 4380 61446
rect 4436 61444 4460 61446
rect 4516 61444 4522 61446
rect 4214 61435 4522 61444
rect 21100 61402 21128 61746
rect 34934 61500 35242 61509
rect 34934 61498 34940 61500
rect 34996 61498 35020 61500
rect 35076 61498 35100 61500
rect 35156 61498 35180 61500
rect 35236 61498 35242 61500
rect 34996 61446 34998 61498
rect 35178 61446 35180 61498
rect 34934 61444 34940 61446
rect 34996 61444 35020 61446
rect 35076 61444 35100 61446
rect 35156 61444 35180 61446
rect 35236 61444 35242 61446
rect 34934 61435 35242 61444
rect 21088 61396 21140 61402
rect 21088 61338 21140 61344
rect 28172 61260 28224 61266
rect 28172 61202 28224 61208
rect 22836 61192 22888 61198
rect 22836 61134 22888 61140
rect 4874 60956 5182 60965
rect 4874 60954 4880 60956
rect 4936 60954 4960 60956
rect 5016 60954 5040 60956
rect 5096 60954 5120 60956
rect 5176 60954 5182 60956
rect 4936 60902 4938 60954
rect 5118 60902 5120 60954
rect 4874 60900 4880 60902
rect 4936 60900 4960 60902
rect 5016 60900 5040 60902
rect 5096 60900 5120 60902
rect 5176 60900 5182 60902
rect 4874 60891 5182 60900
rect 22848 60518 22876 61134
rect 24032 60648 24084 60654
rect 24032 60590 24084 60596
rect 1860 60512 1912 60518
rect 1860 60454 1912 60460
rect 22376 60512 22428 60518
rect 22376 60454 22428 60460
rect 22836 60512 22888 60518
rect 22836 60454 22888 60460
rect 1312 60412 1448 60421
rect 1368 60410 1392 60412
rect 1374 60358 1386 60410
rect 1368 60356 1392 60358
rect 1312 60347 1448 60356
rect 4214 60412 4522 60421
rect 4214 60410 4220 60412
rect 4276 60410 4300 60412
rect 4356 60410 4380 60412
rect 4436 60410 4460 60412
rect 4516 60410 4522 60412
rect 4276 60358 4278 60410
rect 4458 60358 4460 60410
rect 4214 60356 4220 60358
rect 4276 60356 4300 60358
rect 4356 60356 4380 60358
rect 4436 60356 4460 60358
rect 4516 60356 4522 60358
rect 4214 60347 4522 60356
rect 1680 59868 1816 59877
rect 1736 59866 1760 59868
rect 1742 59814 1754 59866
rect 1736 59812 1760 59814
rect 1680 59803 1816 59812
rect 4874 59868 5182 59877
rect 4874 59866 4880 59868
rect 4936 59866 4960 59868
rect 5016 59866 5040 59868
rect 5096 59866 5120 59868
rect 5176 59866 5182 59868
rect 4936 59814 4938 59866
rect 5118 59814 5120 59866
rect 4874 59812 4880 59814
rect 4936 59812 4960 59814
rect 5016 59812 5040 59814
rect 5096 59812 5120 59814
rect 5176 59812 5182 59814
rect 4874 59803 5182 59812
rect 22388 59430 22416 60454
rect 24044 60314 24072 60590
rect 24032 60308 24084 60314
rect 24032 60250 24084 60256
rect 2688 59424 2740 59430
rect 2688 59366 2740 59372
rect 22376 59424 22428 59430
rect 22376 59366 22428 59372
rect 1312 59324 1448 59333
rect 1368 59322 1392 59324
rect 1374 59270 1386 59322
rect 1368 59268 1392 59270
rect 1312 59259 1448 59268
rect 1680 58780 1816 58789
rect 1736 58778 1760 58780
rect 1742 58726 1754 58778
rect 1736 58724 1760 58726
rect 1680 58715 1816 58724
rect 1312 58236 1448 58245
rect 1368 58234 1392 58236
rect 1374 58182 1386 58234
rect 1368 58180 1392 58182
rect 1312 58171 1448 58180
rect 1680 57692 1816 57701
rect 1736 57690 1760 57692
rect 1742 57638 1754 57690
rect 1736 57636 1760 57638
rect 1680 57627 1816 57636
rect 1312 57148 1448 57157
rect 1368 57146 1392 57148
rect 1374 57094 1386 57146
rect 1368 57092 1392 57094
rect 1312 57083 1448 57092
rect 1680 56604 1816 56613
rect 1736 56602 1760 56604
rect 1742 56550 1754 56602
rect 1736 56548 1760 56550
rect 1680 56539 1816 56548
rect 1312 56060 1448 56069
rect 1368 56058 1392 56060
rect 1374 56006 1386 56058
rect 1368 56004 1392 56006
rect 1312 55995 1448 56004
rect 1680 55516 1816 55525
rect 1736 55514 1760 55516
rect 1742 55462 1754 55514
rect 1736 55460 1760 55462
rect 1680 55451 1816 55460
rect 1312 54972 1448 54981
rect 1368 54970 1392 54972
rect 1374 54918 1386 54970
rect 1368 54916 1392 54918
rect 1312 54907 1448 54916
rect 1680 54428 1816 54437
rect 1736 54426 1760 54428
rect 1742 54374 1754 54426
rect 1736 54372 1760 54374
rect 1680 54363 1816 54372
rect 1312 53884 1448 53893
rect 1368 53882 1392 53884
rect 1374 53830 1386 53882
rect 1368 53828 1392 53830
rect 1312 53819 1448 53828
rect 1680 53340 1816 53349
rect 1736 53338 1760 53340
rect 1742 53286 1754 53338
rect 1736 53284 1760 53286
rect 1680 53275 1816 53284
rect 1312 52796 1448 52805
rect 1368 52794 1392 52796
rect 1374 52742 1386 52794
rect 1368 52740 1392 52742
rect 1312 52731 1448 52740
rect 1680 52252 1816 52261
rect 1736 52250 1760 52252
rect 1742 52198 1754 52250
rect 1736 52196 1760 52198
rect 1680 52187 1816 52196
rect 1312 51708 1448 51717
rect 1368 51706 1392 51708
rect 1374 51654 1386 51706
rect 1368 51652 1392 51654
rect 1312 51643 1448 51652
rect 1680 51164 1816 51173
rect 1736 51162 1760 51164
rect 1742 51110 1754 51162
rect 1736 51108 1760 51110
rect 1680 51099 1816 51108
rect 1312 50620 1448 50629
rect 1368 50618 1392 50620
rect 1374 50566 1386 50618
rect 1368 50564 1392 50566
rect 1312 50555 1448 50564
rect 1680 50076 1816 50085
rect 1736 50074 1760 50076
rect 1742 50022 1754 50074
rect 1736 50020 1760 50022
rect 1680 50011 1816 50020
rect 1312 49532 1448 49541
rect 1368 49530 1392 49532
rect 1374 49478 1386 49530
rect 1368 49476 1392 49478
rect 1312 49467 1448 49476
rect 1680 48988 1816 48997
rect 1736 48986 1760 48988
rect 1742 48934 1754 48986
rect 1736 48932 1760 48934
rect 1680 48923 1816 48932
rect 1312 48444 1448 48453
rect 1368 48442 1392 48444
rect 1374 48390 1386 48442
rect 1368 48388 1392 48390
rect 1312 48379 1448 48388
rect 1680 47900 1816 47909
rect 1736 47898 1760 47900
rect 1742 47846 1754 47898
rect 1736 47844 1760 47846
rect 1680 47835 1816 47844
rect 1312 47356 1448 47365
rect 1368 47354 1392 47356
rect 1374 47302 1386 47354
rect 1368 47300 1392 47302
rect 1312 47291 1448 47300
rect 1680 46812 1816 46821
rect 1736 46810 1760 46812
rect 1742 46758 1754 46810
rect 1736 46756 1760 46758
rect 1680 46747 1816 46756
rect 1312 46268 1448 46277
rect 1368 46266 1392 46268
rect 1374 46214 1386 46266
rect 1368 46212 1392 46214
rect 1312 46203 1448 46212
rect 1680 45724 1816 45733
rect 1736 45722 1760 45724
rect 1742 45670 1754 45722
rect 1736 45668 1760 45670
rect 1680 45659 1816 45668
rect 1312 45180 1448 45189
rect 1368 45178 1392 45180
rect 1374 45126 1386 45178
rect 1368 45124 1392 45126
rect 1312 45115 1448 45124
rect 1680 44636 1816 44645
rect 1736 44634 1760 44636
rect 1742 44582 1754 44634
rect 1736 44580 1760 44582
rect 1680 44571 1816 44580
rect 1312 44092 1448 44101
rect 1368 44090 1392 44092
rect 1374 44038 1386 44090
rect 1368 44036 1392 44038
rect 1312 44027 1448 44036
rect 1680 43548 1816 43557
rect 1736 43546 1760 43548
rect 1742 43494 1754 43546
rect 1736 43492 1760 43494
rect 1680 43483 1816 43492
rect 1312 43004 1448 43013
rect 1368 43002 1392 43004
rect 1374 42950 1386 43002
rect 1368 42948 1392 42950
rect 1312 42939 1448 42948
rect 1680 42460 1816 42469
rect 1736 42458 1760 42460
rect 1742 42406 1754 42458
rect 1736 42404 1760 42406
rect 1680 42395 1816 42404
rect 1312 41916 1448 41925
rect 1368 41914 1392 41916
rect 1374 41862 1386 41914
rect 1368 41860 1392 41862
rect 1312 41851 1448 41860
rect 1680 41372 1816 41381
rect 1736 41370 1760 41372
rect 1742 41318 1754 41370
rect 1736 41316 1760 41318
rect 1680 41307 1816 41316
rect 1312 40828 1448 40837
rect 1368 40826 1392 40828
rect 1374 40774 1386 40826
rect 1368 40772 1392 40774
rect 1312 40763 1448 40772
rect 1680 40284 1816 40293
rect 1736 40282 1760 40284
rect 1742 40230 1754 40282
rect 1736 40228 1760 40230
rect 1680 40219 1816 40228
rect 1312 39740 1448 39749
rect 1368 39738 1392 39740
rect 1374 39686 1386 39738
rect 1368 39684 1392 39686
rect 1312 39675 1448 39684
rect 1680 39196 1816 39205
rect 1736 39194 1760 39196
rect 1742 39142 1754 39194
rect 1736 39140 1760 39142
rect 1680 39131 1816 39140
rect 1312 38652 1448 38661
rect 1368 38650 1392 38652
rect 1374 38598 1386 38650
rect 1368 38596 1392 38598
rect 1312 38587 1448 38596
rect 1680 38108 1816 38117
rect 1736 38106 1760 38108
rect 1742 38054 1754 38106
rect 1736 38052 1760 38054
rect 1680 38043 1816 38052
rect 1312 37564 1448 37573
rect 1368 37562 1392 37564
rect 1374 37510 1386 37562
rect 1368 37508 1392 37510
rect 1312 37499 1448 37508
rect 1680 37020 1816 37029
rect 1736 37018 1760 37020
rect 1742 36966 1754 37018
rect 1736 36964 1760 36966
rect 1680 36955 1816 36964
rect 1312 36476 1448 36485
rect 1368 36474 1392 36476
rect 1374 36422 1386 36474
rect 1368 36420 1392 36422
rect 1312 36411 1448 36420
rect 1680 35932 1816 35941
rect 1736 35930 1760 35932
rect 1742 35878 1754 35930
rect 1736 35876 1760 35878
rect 1680 35867 1816 35876
rect 1312 35388 1448 35397
rect 1368 35386 1392 35388
rect 1374 35334 1386 35386
rect 1368 35332 1392 35334
rect 1312 35323 1448 35332
rect 1680 34844 1816 34853
rect 1736 34842 1760 34844
rect 1742 34790 1754 34842
rect 1736 34788 1760 34790
rect 1680 34779 1816 34788
rect 1312 34300 1448 34309
rect 1368 34298 1392 34300
rect 1374 34246 1386 34298
rect 1368 34244 1392 34246
rect 1312 34235 1448 34244
rect 1680 33756 1816 33765
rect 1736 33754 1760 33756
rect 1742 33702 1754 33754
rect 1736 33700 1760 33702
rect 1680 33691 1816 33700
rect 1312 33212 1448 33221
rect 1368 33210 1392 33212
rect 1374 33158 1386 33210
rect 1368 33156 1392 33158
rect 1312 33147 1448 33156
rect 1680 32668 1816 32677
rect 1736 32666 1760 32668
rect 1742 32614 1754 32666
rect 1736 32612 1760 32614
rect 1680 32603 1816 32612
rect 1312 32124 1448 32133
rect 1368 32122 1392 32124
rect 1374 32070 1386 32122
rect 1368 32068 1392 32070
rect 1312 32059 1448 32068
rect 1680 31580 1816 31589
rect 1736 31578 1760 31580
rect 1742 31526 1754 31578
rect 1736 31524 1760 31526
rect 1680 31515 1816 31524
rect 1312 31036 1448 31045
rect 1368 31034 1392 31036
rect 1374 30982 1386 31034
rect 1368 30980 1392 30982
rect 1312 30971 1448 30980
rect 1680 30492 1816 30501
rect 1736 30490 1760 30492
rect 1742 30438 1754 30490
rect 1736 30436 1760 30438
rect 1680 30427 1816 30436
rect 1312 29948 1448 29957
rect 1368 29946 1392 29948
rect 1374 29894 1386 29946
rect 1368 29892 1392 29894
rect 1312 29883 1448 29892
rect 1680 29404 1816 29413
rect 1736 29402 1760 29404
rect 1742 29350 1754 29402
rect 1736 29348 1760 29350
rect 1680 29339 1816 29348
rect 1312 28860 1448 28869
rect 1368 28858 1392 28860
rect 1374 28806 1386 28858
rect 1368 28804 1392 28806
rect 1312 28795 1448 28804
rect 1680 28316 1816 28325
rect 1736 28314 1760 28316
rect 1742 28262 1754 28314
rect 1736 28260 1760 28262
rect 1680 28251 1816 28260
rect 1312 27772 1448 27781
rect 1368 27770 1392 27772
rect 1374 27718 1386 27770
rect 1368 27716 1392 27718
rect 1312 27707 1448 27716
rect 1680 27228 1816 27237
rect 1736 27226 1760 27228
rect 1742 27174 1754 27226
rect 1736 27172 1760 27174
rect 1680 27163 1816 27172
rect 1312 26684 1448 26693
rect 1368 26682 1392 26684
rect 1374 26630 1386 26682
rect 1368 26628 1392 26630
rect 1312 26619 1448 26628
rect 1680 26140 1816 26149
rect 1736 26138 1760 26140
rect 1742 26086 1754 26138
rect 1736 26084 1760 26086
rect 1680 26075 1816 26084
rect 1312 25596 1448 25605
rect 1368 25594 1392 25596
rect 1374 25542 1386 25594
rect 1368 25540 1392 25542
rect 1312 25531 1448 25540
rect 1680 25052 1816 25061
rect 1736 25050 1760 25052
rect 1742 24998 1754 25050
rect 1736 24996 1760 24998
rect 1680 24987 1816 24996
rect 1312 24508 1448 24517
rect 1368 24506 1392 24508
rect 1374 24454 1386 24506
rect 1368 24452 1392 24454
rect 1312 24443 1448 24452
rect 1680 23964 1816 23973
rect 1736 23962 1760 23964
rect 1742 23910 1754 23962
rect 1736 23908 1760 23910
rect 1680 23899 1816 23908
rect 1312 23420 1448 23429
rect 1368 23418 1392 23420
rect 1374 23366 1386 23418
rect 1368 23364 1392 23366
rect 1312 23355 1448 23364
rect 1680 22876 1816 22885
rect 1736 22874 1760 22876
rect 1742 22822 1754 22874
rect 1736 22820 1760 22822
rect 1680 22811 1816 22820
rect 1312 22332 1448 22341
rect 1368 22330 1392 22332
rect 1374 22278 1386 22330
rect 1368 22276 1392 22278
rect 1312 22267 1448 22276
rect 1680 21788 1816 21797
rect 1736 21786 1760 21788
rect 1742 21734 1754 21786
rect 1736 21732 1760 21734
rect 1680 21723 1816 21732
rect 1312 21244 1448 21253
rect 1368 21242 1392 21244
rect 1374 21190 1386 21242
rect 1368 21188 1392 21190
rect 1312 21179 1448 21188
rect 1680 20700 1816 20709
rect 1736 20698 1760 20700
rect 1742 20646 1754 20698
rect 1736 20644 1760 20646
rect 1680 20635 1816 20644
rect 1312 20156 1448 20165
rect 1368 20154 1392 20156
rect 1374 20102 1386 20154
rect 1368 20100 1392 20102
rect 1312 20091 1448 20100
rect 1680 19612 1816 19621
rect 1736 19610 1760 19612
rect 1742 19558 1754 19610
rect 1736 19556 1760 19558
rect 1680 19547 1816 19556
rect 1312 19068 1448 19077
rect 1368 19066 1392 19068
rect 1374 19014 1386 19066
rect 1368 19012 1392 19014
rect 1312 19003 1448 19012
rect 1680 18524 1816 18533
rect 1736 18522 1760 18524
rect 1742 18470 1754 18522
rect 1736 18468 1760 18470
rect 1680 18459 1816 18468
rect 1312 17980 1448 17989
rect 1368 17978 1392 17980
rect 1374 17926 1386 17978
rect 1368 17924 1392 17926
rect 1312 17915 1448 17924
rect 1680 17436 1816 17445
rect 1736 17434 1760 17436
rect 1742 17382 1754 17434
rect 1736 17380 1760 17382
rect 1680 17371 1816 17380
rect 1312 16892 1448 16901
rect 1368 16890 1392 16892
rect 1374 16838 1386 16890
rect 1368 16836 1392 16838
rect 1312 16827 1448 16836
rect 1680 16348 1816 16357
rect 1736 16346 1760 16348
rect 1742 16294 1754 16346
rect 1736 16292 1760 16294
rect 1680 16283 1816 16292
rect 1312 15804 1448 15813
rect 1368 15802 1392 15804
rect 1374 15750 1386 15802
rect 1368 15748 1392 15750
rect 1312 15739 1448 15748
rect 1680 15260 1816 15269
rect 1736 15258 1760 15260
rect 1742 15206 1754 15258
rect 1736 15204 1760 15206
rect 1680 15195 1816 15204
rect 1312 14716 1448 14725
rect 1368 14714 1392 14716
rect 1374 14662 1386 14714
rect 1368 14660 1392 14662
rect 1312 14651 1448 14660
rect 1680 14172 1816 14181
rect 1736 14170 1760 14172
rect 1742 14118 1754 14170
rect 1736 14116 1760 14118
rect 1680 14107 1816 14116
rect 1312 13628 1448 13637
rect 1368 13626 1392 13628
rect 1374 13574 1386 13626
rect 1368 13572 1392 13574
rect 1312 13563 1448 13572
rect 1680 13084 1816 13093
rect 1736 13082 1760 13084
rect 1742 13030 1754 13082
rect 1736 13028 1760 13030
rect 1680 13019 1816 13028
rect 1312 12540 1448 12549
rect 1368 12538 1392 12540
rect 1374 12486 1386 12538
rect 1368 12484 1392 12486
rect 1312 12475 1448 12484
rect 1680 11996 1816 12005
rect 1736 11994 1760 11996
rect 1742 11942 1754 11994
rect 1736 11940 1760 11942
rect 1680 11931 1816 11940
rect 1312 11452 1448 11461
rect 1368 11450 1392 11452
rect 1374 11398 1386 11450
rect 1368 11396 1392 11398
rect 1312 11387 1448 11396
rect 1680 10908 1816 10917
rect 1736 10906 1760 10908
rect 1742 10854 1754 10906
rect 1736 10852 1760 10854
rect 1680 10843 1816 10852
rect 1312 10364 1448 10373
rect 1368 10362 1392 10364
rect 1374 10310 1386 10362
rect 1368 10308 1392 10310
rect 1312 10299 1448 10308
rect 1680 9820 1816 9829
rect 1736 9818 1760 9820
rect 1742 9766 1754 9818
rect 1736 9764 1760 9766
rect 1680 9755 1816 9764
rect 1312 9276 1448 9285
rect 1368 9274 1392 9276
rect 1374 9222 1386 9274
rect 1368 9220 1392 9222
rect 1312 9211 1448 9220
rect 1680 8732 1816 8741
rect 1736 8730 1760 8732
rect 1742 8678 1754 8730
rect 1736 8676 1760 8678
rect 1680 8667 1816 8676
rect 1312 8188 1448 8197
rect 1368 8186 1392 8188
rect 1374 8134 1386 8186
rect 1368 8132 1392 8134
rect 1312 8123 1448 8132
rect 1680 7644 1816 7653
rect 1736 7642 1760 7644
rect 1742 7590 1754 7642
rect 1736 7588 1760 7590
rect 1680 7579 1816 7588
rect 1312 7100 1448 7109
rect 1368 7098 1392 7100
rect 1374 7046 1386 7098
rect 1368 7044 1392 7046
rect 1312 7035 1448 7044
rect 1680 6556 1816 6565
rect 1736 6554 1760 6556
rect 1742 6502 1754 6554
rect 1736 6500 1760 6502
rect 1680 6491 1816 6500
rect 1312 6012 1448 6021
rect 1368 6010 1392 6012
rect 1374 5958 1386 6010
rect 1368 5956 1392 5958
rect 1312 5947 1448 5956
rect 1680 5468 1816 5477
rect 1736 5466 1760 5468
rect 1742 5414 1754 5466
rect 1736 5412 1760 5414
rect 1680 5403 1816 5412
rect 1312 4924 1448 4933
rect 1368 4922 1392 4924
rect 1374 4870 1386 4922
rect 1368 4868 1392 4870
rect 1312 4859 1448 4868
rect 1680 4380 1816 4389
rect 1736 4378 1760 4380
rect 1742 4326 1754 4378
rect 1736 4324 1760 4326
rect 1680 4315 1816 4324
rect 2700 3913 2728 59366
rect 28184 57905 28212 61202
rect 28816 61056 28868 61062
rect 28816 60998 28868 61004
rect 28828 60722 28856 60998
rect 35594 60956 35902 60965
rect 35594 60954 35600 60956
rect 35656 60954 35680 60956
rect 35736 60954 35760 60956
rect 35816 60954 35840 60956
rect 35896 60954 35902 60956
rect 35656 60902 35658 60954
rect 35838 60902 35840 60954
rect 35594 60900 35600 60902
rect 35656 60900 35680 60902
rect 35736 60900 35760 60902
rect 35816 60900 35840 60902
rect 35896 60900 35902 60902
rect 35594 60891 35902 60900
rect 46676 60722 46704 74802
rect 49436 60790 49464 76978
rect 49620 76634 49648 77007
rect 49608 76628 49660 76634
rect 49608 76570 49660 76576
rect 49988 75002 50016 77318
rect 51092 75002 51120 77386
rect 51184 77178 51212 101390
rect 53116 77722 53144 101390
rect 55140 77722 55168 101390
rect 57348 77722 57376 101390
rect 59188 77722 59216 101390
rect 66314 101212 66622 101221
rect 66314 101210 66320 101212
rect 66376 101210 66400 101212
rect 66456 101210 66480 101212
rect 66536 101210 66560 101212
rect 66616 101210 66622 101212
rect 66376 101158 66378 101210
rect 66558 101158 66560 101210
rect 66314 101156 66320 101158
rect 66376 101156 66400 101158
rect 66456 101156 66480 101158
rect 66536 101156 66560 101158
rect 66616 101156 66622 101158
rect 66314 101147 66622 101156
rect 97034 101212 97342 101221
rect 97034 101210 97040 101212
rect 97096 101210 97120 101212
rect 97176 101210 97200 101212
rect 97256 101210 97280 101212
rect 97336 101210 97342 101212
rect 97096 101158 97098 101210
rect 97278 101158 97280 101210
rect 97034 101156 97040 101158
rect 97096 101156 97120 101158
rect 97176 101156 97200 101158
rect 97256 101156 97280 101158
rect 97336 101156 97342 101158
rect 97034 101147 97342 101156
rect 65654 100668 65962 100677
rect 65654 100666 65660 100668
rect 65716 100666 65740 100668
rect 65796 100666 65820 100668
rect 65876 100666 65900 100668
rect 65956 100666 65962 100668
rect 65716 100614 65718 100666
rect 65898 100614 65900 100666
rect 65654 100612 65660 100614
rect 65716 100612 65740 100614
rect 65796 100612 65820 100614
rect 65876 100612 65900 100614
rect 65956 100612 65962 100614
rect 65654 100603 65962 100612
rect 96374 100668 96682 100677
rect 96374 100666 96380 100668
rect 96436 100666 96460 100668
rect 96516 100666 96540 100668
rect 96596 100666 96620 100668
rect 96676 100666 96682 100668
rect 96436 100614 96438 100666
rect 96618 100614 96620 100666
rect 96374 100612 96380 100614
rect 96436 100612 96460 100614
rect 96516 100612 96540 100614
rect 96596 100612 96620 100614
rect 96676 100612 96682 100614
rect 96374 100603 96682 100612
rect 66314 100124 66622 100133
rect 66314 100122 66320 100124
rect 66376 100122 66400 100124
rect 66456 100122 66480 100124
rect 66536 100122 66560 100124
rect 66616 100122 66622 100124
rect 66376 100070 66378 100122
rect 66558 100070 66560 100122
rect 66314 100068 66320 100070
rect 66376 100068 66400 100070
rect 66456 100068 66480 100070
rect 66536 100068 66560 100070
rect 66616 100068 66622 100070
rect 66314 100059 66622 100068
rect 97034 100124 97342 100133
rect 97034 100122 97040 100124
rect 97096 100122 97120 100124
rect 97176 100122 97200 100124
rect 97256 100122 97280 100124
rect 97336 100122 97342 100124
rect 97096 100070 97098 100122
rect 97278 100070 97280 100122
rect 97034 100068 97040 100070
rect 97096 100068 97120 100070
rect 97176 100068 97200 100070
rect 97256 100068 97280 100070
rect 97336 100068 97342 100070
rect 97034 100059 97342 100068
rect 65654 99580 65962 99589
rect 65654 99578 65660 99580
rect 65716 99578 65740 99580
rect 65796 99578 65820 99580
rect 65876 99578 65900 99580
rect 65956 99578 65962 99580
rect 65716 99526 65718 99578
rect 65898 99526 65900 99578
rect 65654 99524 65660 99526
rect 65716 99524 65740 99526
rect 65796 99524 65820 99526
rect 65876 99524 65900 99526
rect 65956 99524 65962 99526
rect 65654 99515 65962 99524
rect 96374 99580 96682 99589
rect 96374 99578 96380 99580
rect 96436 99578 96460 99580
rect 96516 99578 96540 99580
rect 96596 99578 96620 99580
rect 96676 99578 96682 99580
rect 96436 99526 96438 99578
rect 96618 99526 96620 99578
rect 96374 99524 96380 99526
rect 96436 99524 96460 99526
rect 96516 99524 96540 99526
rect 96596 99524 96620 99526
rect 96676 99524 96682 99526
rect 96374 99515 96682 99524
rect 66314 99036 66622 99045
rect 66314 99034 66320 99036
rect 66376 99034 66400 99036
rect 66456 99034 66480 99036
rect 66536 99034 66560 99036
rect 66616 99034 66622 99036
rect 66376 98982 66378 99034
rect 66558 98982 66560 99034
rect 66314 98980 66320 98982
rect 66376 98980 66400 98982
rect 66456 98980 66480 98982
rect 66536 98980 66560 98982
rect 66616 98980 66622 98982
rect 66314 98971 66622 98980
rect 97034 99036 97342 99045
rect 97034 99034 97040 99036
rect 97096 99034 97120 99036
rect 97176 99034 97200 99036
rect 97256 99034 97280 99036
rect 97336 99034 97342 99036
rect 97096 98982 97098 99034
rect 97278 98982 97280 99034
rect 97034 98980 97040 98982
rect 97096 98980 97120 98982
rect 97176 98980 97200 98982
rect 97256 98980 97280 98982
rect 97336 98980 97342 98982
rect 97034 98971 97342 98980
rect 65654 98492 65962 98501
rect 65654 98490 65660 98492
rect 65716 98490 65740 98492
rect 65796 98490 65820 98492
rect 65876 98490 65900 98492
rect 65956 98490 65962 98492
rect 65716 98438 65718 98490
rect 65898 98438 65900 98490
rect 65654 98436 65660 98438
rect 65716 98436 65740 98438
rect 65796 98436 65820 98438
rect 65876 98436 65900 98438
rect 65956 98436 65962 98438
rect 65654 98427 65962 98436
rect 96374 98492 96682 98501
rect 96374 98490 96380 98492
rect 96436 98490 96460 98492
rect 96516 98490 96540 98492
rect 96596 98490 96620 98492
rect 96676 98490 96682 98492
rect 96436 98438 96438 98490
rect 96618 98438 96620 98490
rect 96374 98436 96380 98438
rect 96436 98436 96460 98438
rect 96516 98436 96540 98438
rect 96596 98436 96620 98438
rect 96676 98436 96682 98438
rect 96374 98427 96682 98436
rect 66314 97948 66622 97957
rect 66314 97946 66320 97948
rect 66376 97946 66400 97948
rect 66456 97946 66480 97948
rect 66536 97946 66560 97948
rect 66616 97946 66622 97948
rect 66376 97894 66378 97946
rect 66558 97894 66560 97946
rect 66314 97892 66320 97894
rect 66376 97892 66400 97894
rect 66456 97892 66480 97894
rect 66536 97892 66560 97894
rect 66616 97892 66622 97894
rect 66314 97883 66622 97892
rect 97034 97948 97342 97957
rect 97034 97946 97040 97948
rect 97096 97946 97120 97948
rect 97176 97946 97200 97948
rect 97256 97946 97280 97948
rect 97336 97946 97342 97948
rect 97096 97894 97098 97946
rect 97278 97894 97280 97946
rect 97034 97892 97040 97894
rect 97096 97892 97120 97894
rect 97176 97892 97200 97894
rect 97256 97892 97280 97894
rect 97336 97892 97342 97894
rect 97034 97883 97342 97892
rect 65654 97404 65962 97413
rect 65654 97402 65660 97404
rect 65716 97402 65740 97404
rect 65796 97402 65820 97404
rect 65876 97402 65900 97404
rect 65956 97402 65962 97404
rect 65716 97350 65718 97402
rect 65898 97350 65900 97402
rect 65654 97348 65660 97350
rect 65716 97348 65740 97350
rect 65796 97348 65820 97350
rect 65876 97348 65900 97350
rect 65956 97348 65962 97350
rect 65654 97339 65962 97348
rect 96374 97404 96682 97413
rect 96374 97402 96380 97404
rect 96436 97402 96460 97404
rect 96516 97402 96540 97404
rect 96596 97402 96620 97404
rect 96676 97402 96682 97404
rect 96436 97350 96438 97402
rect 96618 97350 96620 97402
rect 96374 97348 96380 97350
rect 96436 97348 96460 97350
rect 96516 97348 96540 97350
rect 96596 97348 96620 97350
rect 96676 97348 96682 97350
rect 96374 97339 96682 97348
rect 66314 96860 66622 96869
rect 66314 96858 66320 96860
rect 66376 96858 66400 96860
rect 66456 96858 66480 96860
rect 66536 96858 66560 96860
rect 66616 96858 66622 96860
rect 66376 96806 66378 96858
rect 66558 96806 66560 96858
rect 66314 96804 66320 96806
rect 66376 96804 66400 96806
rect 66456 96804 66480 96806
rect 66536 96804 66560 96806
rect 66616 96804 66622 96806
rect 66314 96795 66622 96804
rect 97034 96860 97342 96869
rect 97034 96858 97040 96860
rect 97096 96858 97120 96860
rect 97176 96858 97200 96860
rect 97256 96858 97280 96860
rect 97336 96858 97342 96860
rect 97096 96806 97098 96858
rect 97278 96806 97280 96858
rect 97034 96804 97040 96806
rect 97096 96804 97120 96806
rect 97176 96804 97200 96806
rect 97256 96804 97280 96806
rect 97336 96804 97342 96806
rect 97034 96795 97342 96804
rect 65654 96316 65962 96325
rect 65654 96314 65660 96316
rect 65716 96314 65740 96316
rect 65796 96314 65820 96316
rect 65876 96314 65900 96316
rect 65956 96314 65962 96316
rect 65716 96262 65718 96314
rect 65898 96262 65900 96314
rect 65654 96260 65660 96262
rect 65716 96260 65740 96262
rect 65796 96260 65820 96262
rect 65876 96260 65900 96262
rect 65956 96260 65962 96262
rect 65654 96251 65962 96260
rect 96374 96316 96682 96325
rect 96374 96314 96380 96316
rect 96436 96314 96460 96316
rect 96516 96314 96540 96316
rect 96596 96314 96620 96316
rect 96676 96314 96682 96316
rect 96436 96262 96438 96314
rect 96618 96262 96620 96314
rect 96374 96260 96380 96262
rect 96436 96260 96460 96262
rect 96516 96260 96540 96262
rect 96596 96260 96620 96262
rect 96676 96260 96682 96262
rect 96374 96251 96682 96260
rect 66314 95772 66622 95781
rect 66314 95770 66320 95772
rect 66376 95770 66400 95772
rect 66456 95770 66480 95772
rect 66536 95770 66560 95772
rect 66616 95770 66622 95772
rect 66376 95718 66378 95770
rect 66558 95718 66560 95770
rect 66314 95716 66320 95718
rect 66376 95716 66400 95718
rect 66456 95716 66480 95718
rect 66536 95716 66560 95718
rect 66616 95716 66622 95718
rect 66314 95707 66622 95716
rect 97034 95772 97342 95781
rect 97034 95770 97040 95772
rect 97096 95770 97120 95772
rect 97176 95770 97200 95772
rect 97256 95770 97280 95772
rect 97336 95770 97342 95772
rect 97096 95718 97098 95770
rect 97278 95718 97280 95770
rect 97034 95716 97040 95718
rect 97096 95716 97120 95718
rect 97176 95716 97200 95718
rect 97256 95716 97280 95718
rect 97336 95716 97342 95718
rect 97034 95707 97342 95716
rect 65654 95228 65962 95237
rect 65654 95226 65660 95228
rect 65716 95226 65740 95228
rect 65796 95226 65820 95228
rect 65876 95226 65900 95228
rect 65956 95226 65962 95228
rect 65716 95174 65718 95226
rect 65898 95174 65900 95226
rect 65654 95172 65660 95174
rect 65716 95172 65740 95174
rect 65796 95172 65820 95174
rect 65876 95172 65900 95174
rect 65956 95172 65962 95174
rect 65654 95163 65962 95172
rect 96374 95228 96682 95237
rect 96374 95226 96380 95228
rect 96436 95226 96460 95228
rect 96516 95226 96540 95228
rect 96596 95226 96620 95228
rect 96676 95226 96682 95228
rect 96436 95174 96438 95226
rect 96618 95174 96620 95226
rect 96374 95172 96380 95174
rect 96436 95172 96460 95174
rect 96516 95172 96540 95174
rect 96596 95172 96620 95174
rect 96676 95172 96682 95174
rect 96374 95163 96682 95172
rect 66314 94684 66622 94693
rect 66314 94682 66320 94684
rect 66376 94682 66400 94684
rect 66456 94682 66480 94684
rect 66536 94682 66560 94684
rect 66616 94682 66622 94684
rect 66376 94630 66378 94682
rect 66558 94630 66560 94682
rect 66314 94628 66320 94630
rect 66376 94628 66400 94630
rect 66456 94628 66480 94630
rect 66536 94628 66560 94630
rect 66616 94628 66622 94630
rect 66314 94619 66622 94628
rect 97034 94684 97342 94693
rect 97034 94682 97040 94684
rect 97096 94682 97120 94684
rect 97176 94682 97200 94684
rect 97256 94682 97280 94684
rect 97336 94682 97342 94684
rect 97096 94630 97098 94682
rect 97278 94630 97280 94682
rect 97034 94628 97040 94630
rect 97096 94628 97120 94630
rect 97176 94628 97200 94630
rect 97256 94628 97280 94630
rect 97336 94628 97342 94630
rect 97034 94619 97342 94628
rect 65654 94140 65962 94149
rect 65654 94138 65660 94140
rect 65716 94138 65740 94140
rect 65796 94138 65820 94140
rect 65876 94138 65900 94140
rect 65956 94138 65962 94140
rect 65716 94086 65718 94138
rect 65898 94086 65900 94138
rect 65654 94084 65660 94086
rect 65716 94084 65740 94086
rect 65796 94084 65820 94086
rect 65876 94084 65900 94086
rect 65956 94084 65962 94086
rect 65654 94075 65962 94084
rect 96374 94140 96682 94149
rect 96374 94138 96380 94140
rect 96436 94138 96460 94140
rect 96516 94138 96540 94140
rect 96596 94138 96620 94140
rect 96676 94138 96682 94140
rect 96436 94086 96438 94138
rect 96618 94086 96620 94138
rect 96374 94084 96380 94086
rect 96436 94084 96460 94086
rect 96516 94084 96540 94086
rect 96596 94084 96620 94086
rect 96676 94084 96682 94086
rect 96374 94075 96682 94084
rect 66314 93596 66622 93605
rect 66314 93594 66320 93596
rect 66376 93594 66400 93596
rect 66456 93594 66480 93596
rect 66536 93594 66560 93596
rect 66616 93594 66622 93596
rect 66376 93542 66378 93594
rect 66558 93542 66560 93594
rect 66314 93540 66320 93542
rect 66376 93540 66400 93542
rect 66456 93540 66480 93542
rect 66536 93540 66560 93542
rect 66616 93540 66622 93542
rect 66314 93531 66622 93540
rect 97034 93596 97342 93605
rect 97034 93594 97040 93596
rect 97096 93594 97120 93596
rect 97176 93594 97200 93596
rect 97256 93594 97280 93596
rect 97336 93594 97342 93596
rect 97096 93542 97098 93594
rect 97278 93542 97280 93594
rect 97034 93540 97040 93542
rect 97096 93540 97120 93542
rect 97176 93540 97200 93542
rect 97256 93540 97280 93542
rect 97336 93540 97342 93542
rect 97034 93531 97342 93540
rect 65654 93052 65962 93061
rect 65654 93050 65660 93052
rect 65716 93050 65740 93052
rect 65796 93050 65820 93052
rect 65876 93050 65900 93052
rect 65956 93050 65962 93052
rect 65716 92998 65718 93050
rect 65898 92998 65900 93050
rect 65654 92996 65660 92998
rect 65716 92996 65740 92998
rect 65796 92996 65820 92998
rect 65876 92996 65900 92998
rect 65956 92996 65962 92998
rect 65654 92987 65962 92996
rect 96374 93052 96682 93061
rect 96374 93050 96380 93052
rect 96436 93050 96460 93052
rect 96516 93050 96540 93052
rect 96596 93050 96620 93052
rect 96676 93050 96682 93052
rect 96436 92998 96438 93050
rect 96618 92998 96620 93050
rect 96374 92996 96380 92998
rect 96436 92996 96460 92998
rect 96516 92996 96540 92998
rect 96596 92996 96620 92998
rect 96676 92996 96682 92998
rect 96374 92987 96682 92996
rect 66314 92508 66622 92517
rect 66314 92506 66320 92508
rect 66376 92506 66400 92508
rect 66456 92506 66480 92508
rect 66536 92506 66560 92508
rect 66616 92506 66622 92508
rect 66376 92454 66378 92506
rect 66558 92454 66560 92506
rect 66314 92452 66320 92454
rect 66376 92452 66400 92454
rect 66456 92452 66480 92454
rect 66536 92452 66560 92454
rect 66616 92452 66622 92454
rect 66314 92443 66622 92452
rect 97034 92508 97342 92517
rect 97034 92506 97040 92508
rect 97096 92506 97120 92508
rect 97176 92506 97200 92508
rect 97256 92506 97280 92508
rect 97336 92506 97342 92508
rect 97096 92454 97098 92506
rect 97278 92454 97280 92506
rect 97034 92452 97040 92454
rect 97096 92452 97120 92454
rect 97176 92452 97200 92454
rect 97256 92452 97280 92454
rect 97336 92452 97342 92454
rect 97034 92443 97342 92452
rect 65654 91964 65962 91973
rect 65654 91962 65660 91964
rect 65716 91962 65740 91964
rect 65796 91962 65820 91964
rect 65876 91962 65900 91964
rect 65956 91962 65962 91964
rect 65716 91910 65718 91962
rect 65898 91910 65900 91962
rect 65654 91908 65660 91910
rect 65716 91908 65740 91910
rect 65796 91908 65820 91910
rect 65876 91908 65900 91910
rect 65956 91908 65962 91910
rect 65654 91899 65962 91908
rect 96374 91964 96682 91973
rect 96374 91962 96380 91964
rect 96436 91962 96460 91964
rect 96516 91962 96540 91964
rect 96596 91962 96620 91964
rect 96676 91962 96682 91964
rect 96436 91910 96438 91962
rect 96618 91910 96620 91962
rect 96374 91908 96380 91910
rect 96436 91908 96460 91910
rect 96516 91908 96540 91910
rect 96596 91908 96620 91910
rect 96676 91908 96682 91910
rect 96374 91899 96682 91908
rect 66314 91420 66622 91429
rect 66314 91418 66320 91420
rect 66376 91418 66400 91420
rect 66456 91418 66480 91420
rect 66536 91418 66560 91420
rect 66616 91418 66622 91420
rect 66376 91366 66378 91418
rect 66558 91366 66560 91418
rect 66314 91364 66320 91366
rect 66376 91364 66400 91366
rect 66456 91364 66480 91366
rect 66536 91364 66560 91366
rect 66616 91364 66622 91366
rect 66314 91355 66622 91364
rect 97034 91420 97342 91429
rect 97034 91418 97040 91420
rect 97096 91418 97120 91420
rect 97176 91418 97200 91420
rect 97256 91418 97280 91420
rect 97336 91418 97342 91420
rect 97096 91366 97098 91418
rect 97278 91366 97280 91418
rect 97034 91364 97040 91366
rect 97096 91364 97120 91366
rect 97176 91364 97200 91366
rect 97256 91364 97280 91366
rect 97336 91364 97342 91366
rect 97034 91355 97342 91364
rect 65654 90876 65962 90885
rect 65654 90874 65660 90876
rect 65716 90874 65740 90876
rect 65796 90874 65820 90876
rect 65876 90874 65900 90876
rect 65956 90874 65962 90876
rect 65716 90822 65718 90874
rect 65898 90822 65900 90874
rect 65654 90820 65660 90822
rect 65716 90820 65740 90822
rect 65796 90820 65820 90822
rect 65876 90820 65900 90822
rect 65956 90820 65962 90822
rect 65654 90811 65962 90820
rect 96374 90876 96682 90885
rect 96374 90874 96380 90876
rect 96436 90874 96460 90876
rect 96516 90874 96540 90876
rect 96596 90874 96620 90876
rect 96676 90874 96682 90876
rect 96436 90822 96438 90874
rect 96618 90822 96620 90874
rect 96374 90820 96380 90822
rect 96436 90820 96460 90822
rect 96516 90820 96540 90822
rect 96596 90820 96620 90822
rect 96676 90820 96682 90822
rect 96374 90811 96682 90820
rect 66314 90332 66622 90341
rect 66314 90330 66320 90332
rect 66376 90330 66400 90332
rect 66456 90330 66480 90332
rect 66536 90330 66560 90332
rect 66616 90330 66622 90332
rect 66376 90278 66378 90330
rect 66558 90278 66560 90330
rect 66314 90276 66320 90278
rect 66376 90276 66400 90278
rect 66456 90276 66480 90278
rect 66536 90276 66560 90278
rect 66616 90276 66622 90278
rect 66314 90267 66622 90276
rect 97034 90332 97342 90341
rect 97034 90330 97040 90332
rect 97096 90330 97120 90332
rect 97176 90330 97200 90332
rect 97256 90330 97280 90332
rect 97336 90330 97342 90332
rect 97096 90278 97098 90330
rect 97278 90278 97280 90330
rect 97034 90276 97040 90278
rect 97096 90276 97120 90278
rect 97176 90276 97200 90278
rect 97256 90276 97280 90278
rect 97336 90276 97342 90278
rect 97034 90267 97342 90276
rect 65654 89788 65962 89797
rect 65654 89786 65660 89788
rect 65716 89786 65740 89788
rect 65796 89786 65820 89788
rect 65876 89786 65900 89788
rect 65956 89786 65962 89788
rect 65716 89734 65718 89786
rect 65898 89734 65900 89786
rect 65654 89732 65660 89734
rect 65716 89732 65740 89734
rect 65796 89732 65820 89734
rect 65876 89732 65900 89734
rect 65956 89732 65962 89734
rect 65654 89723 65962 89732
rect 96374 89788 96682 89797
rect 96374 89786 96380 89788
rect 96436 89786 96460 89788
rect 96516 89786 96540 89788
rect 96596 89786 96620 89788
rect 96676 89786 96682 89788
rect 96436 89734 96438 89786
rect 96618 89734 96620 89786
rect 96374 89732 96380 89734
rect 96436 89732 96460 89734
rect 96516 89732 96540 89734
rect 96596 89732 96620 89734
rect 96676 89732 96682 89734
rect 96374 89723 96682 89732
rect 66314 89244 66622 89253
rect 66314 89242 66320 89244
rect 66376 89242 66400 89244
rect 66456 89242 66480 89244
rect 66536 89242 66560 89244
rect 66616 89242 66622 89244
rect 66376 89190 66378 89242
rect 66558 89190 66560 89242
rect 66314 89188 66320 89190
rect 66376 89188 66400 89190
rect 66456 89188 66480 89190
rect 66536 89188 66560 89190
rect 66616 89188 66622 89190
rect 66314 89179 66622 89188
rect 97034 89244 97342 89253
rect 97034 89242 97040 89244
rect 97096 89242 97120 89244
rect 97176 89242 97200 89244
rect 97256 89242 97280 89244
rect 97336 89242 97342 89244
rect 97096 89190 97098 89242
rect 97278 89190 97280 89242
rect 97034 89188 97040 89190
rect 97096 89188 97120 89190
rect 97176 89188 97200 89190
rect 97256 89188 97280 89190
rect 97336 89188 97342 89190
rect 97034 89179 97342 89188
rect 65654 88700 65962 88709
rect 65654 88698 65660 88700
rect 65716 88698 65740 88700
rect 65796 88698 65820 88700
rect 65876 88698 65900 88700
rect 65956 88698 65962 88700
rect 65716 88646 65718 88698
rect 65898 88646 65900 88698
rect 65654 88644 65660 88646
rect 65716 88644 65740 88646
rect 65796 88644 65820 88646
rect 65876 88644 65900 88646
rect 65956 88644 65962 88646
rect 65654 88635 65962 88644
rect 96374 88700 96682 88709
rect 96374 88698 96380 88700
rect 96436 88698 96460 88700
rect 96516 88698 96540 88700
rect 96596 88698 96620 88700
rect 96676 88698 96682 88700
rect 96436 88646 96438 88698
rect 96618 88646 96620 88698
rect 96374 88644 96380 88646
rect 96436 88644 96460 88646
rect 96516 88644 96540 88646
rect 96596 88644 96620 88646
rect 96676 88644 96682 88646
rect 96374 88635 96682 88644
rect 66314 88156 66622 88165
rect 66314 88154 66320 88156
rect 66376 88154 66400 88156
rect 66456 88154 66480 88156
rect 66536 88154 66560 88156
rect 66616 88154 66622 88156
rect 66376 88102 66378 88154
rect 66558 88102 66560 88154
rect 66314 88100 66320 88102
rect 66376 88100 66400 88102
rect 66456 88100 66480 88102
rect 66536 88100 66560 88102
rect 66616 88100 66622 88102
rect 66314 88091 66622 88100
rect 97034 88156 97342 88165
rect 97034 88154 97040 88156
rect 97096 88154 97120 88156
rect 97176 88154 97200 88156
rect 97256 88154 97280 88156
rect 97336 88154 97342 88156
rect 97096 88102 97098 88154
rect 97278 88102 97280 88154
rect 97034 88100 97040 88102
rect 97096 88100 97120 88102
rect 97176 88100 97200 88102
rect 97256 88100 97280 88102
rect 97336 88100 97342 88102
rect 97034 88091 97342 88100
rect 65654 87612 65962 87621
rect 65654 87610 65660 87612
rect 65716 87610 65740 87612
rect 65796 87610 65820 87612
rect 65876 87610 65900 87612
rect 65956 87610 65962 87612
rect 65716 87558 65718 87610
rect 65898 87558 65900 87610
rect 65654 87556 65660 87558
rect 65716 87556 65740 87558
rect 65796 87556 65820 87558
rect 65876 87556 65900 87558
rect 65956 87556 65962 87558
rect 65654 87547 65962 87556
rect 96374 87612 96682 87621
rect 96374 87610 96380 87612
rect 96436 87610 96460 87612
rect 96516 87610 96540 87612
rect 96596 87610 96620 87612
rect 96676 87610 96682 87612
rect 96436 87558 96438 87610
rect 96618 87558 96620 87610
rect 96374 87556 96380 87558
rect 96436 87556 96460 87558
rect 96516 87556 96540 87558
rect 96596 87556 96620 87558
rect 96676 87556 96682 87558
rect 96374 87547 96682 87556
rect 66314 87068 66622 87077
rect 66314 87066 66320 87068
rect 66376 87066 66400 87068
rect 66456 87066 66480 87068
rect 66536 87066 66560 87068
rect 66616 87066 66622 87068
rect 66376 87014 66378 87066
rect 66558 87014 66560 87066
rect 66314 87012 66320 87014
rect 66376 87012 66400 87014
rect 66456 87012 66480 87014
rect 66536 87012 66560 87014
rect 66616 87012 66622 87014
rect 66314 87003 66622 87012
rect 97034 87068 97342 87077
rect 97034 87066 97040 87068
rect 97096 87066 97120 87068
rect 97176 87066 97200 87068
rect 97256 87066 97280 87068
rect 97336 87066 97342 87068
rect 97096 87014 97098 87066
rect 97278 87014 97280 87066
rect 97034 87012 97040 87014
rect 97096 87012 97120 87014
rect 97176 87012 97200 87014
rect 97256 87012 97280 87014
rect 97336 87012 97342 87014
rect 97034 87003 97342 87012
rect 65654 86524 65962 86533
rect 65654 86522 65660 86524
rect 65716 86522 65740 86524
rect 65796 86522 65820 86524
rect 65876 86522 65900 86524
rect 65956 86522 65962 86524
rect 65716 86470 65718 86522
rect 65898 86470 65900 86522
rect 65654 86468 65660 86470
rect 65716 86468 65740 86470
rect 65796 86468 65820 86470
rect 65876 86468 65900 86470
rect 65956 86468 65962 86470
rect 65654 86459 65962 86468
rect 96374 86524 96682 86533
rect 96374 86522 96380 86524
rect 96436 86522 96460 86524
rect 96516 86522 96540 86524
rect 96596 86522 96620 86524
rect 96676 86522 96682 86524
rect 96436 86470 96438 86522
rect 96618 86470 96620 86522
rect 96374 86468 96380 86470
rect 96436 86468 96460 86470
rect 96516 86468 96540 86470
rect 96596 86468 96620 86470
rect 96676 86468 96682 86470
rect 96374 86459 96682 86468
rect 66314 85980 66622 85989
rect 66314 85978 66320 85980
rect 66376 85978 66400 85980
rect 66456 85978 66480 85980
rect 66536 85978 66560 85980
rect 66616 85978 66622 85980
rect 66376 85926 66378 85978
rect 66558 85926 66560 85978
rect 66314 85924 66320 85926
rect 66376 85924 66400 85926
rect 66456 85924 66480 85926
rect 66536 85924 66560 85926
rect 66616 85924 66622 85926
rect 66314 85915 66622 85924
rect 97034 85980 97342 85989
rect 97034 85978 97040 85980
rect 97096 85978 97120 85980
rect 97176 85978 97200 85980
rect 97256 85978 97280 85980
rect 97336 85978 97342 85980
rect 97096 85926 97098 85978
rect 97278 85926 97280 85978
rect 97034 85924 97040 85926
rect 97096 85924 97120 85926
rect 97176 85924 97200 85926
rect 97256 85924 97280 85926
rect 97336 85924 97342 85926
rect 97034 85915 97342 85924
rect 65654 85436 65962 85445
rect 65654 85434 65660 85436
rect 65716 85434 65740 85436
rect 65796 85434 65820 85436
rect 65876 85434 65900 85436
rect 65956 85434 65962 85436
rect 65716 85382 65718 85434
rect 65898 85382 65900 85434
rect 65654 85380 65660 85382
rect 65716 85380 65740 85382
rect 65796 85380 65820 85382
rect 65876 85380 65900 85382
rect 65956 85380 65962 85382
rect 65654 85371 65962 85380
rect 96374 85436 96682 85445
rect 96374 85434 96380 85436
rect 96436 85434 96460 85436
rect 96516 85434 96540 85436
rect 96596 85434 96620 85436
rect 96676 85434 96682 85436
rect 96436 85382 96438 85434
rect 96618 85382 96620 85434
rect 96374 85380 96380 85382
rect 96436 85380 96460 85382
rect 96516 85380 96540 85382
rect 96596 85380 96620 85382
rect 96676 85380 96682 85382
rect 96374 85371 96682 85380
rect 66314 84892 66622 84901
rect 66314 84890 66320 84892
rect 66376 84890 66400 84892
rect 66456 84890 66480 84892
rect 66536 84890 66560 84892
rect 66616 84890 66622 84892
rect 66376 84838 66378 84890
rect 66558 84838 66560 84890
rect 66314 84836 66320 84838
rect 66376 84836 66400 84838
rect 66456 84836 66480 84838
rect 66536 84836 66560 84838
rect 66616 84836 66622 84838
rect 66314 84827 66622 84836
rect 97034 84892 97342 84901
rect 97034 84890 97040 84892
rect 97096 84890 97120 84892
rect 97176 84890 97200 84892
rect 97256 84890 97280 84892
rect 97336 84890 97342 84892
rect 97096 84838 97098 84890
rect 97278 84838 97280 84890
rect 97034 84836 97040 84838
rect 97096 84836 97120 84838
rect 97176 84836 97200 84838
rect 97256 84836 97280 84838
rect 97336 84836 97342 84838
rect 97034 84827 97342 84836
rect 65654 84348 65962 84357
rect 65654 84346 65660 84348
rect 65716 84346 65740 84348
rect 65796 84346 65820 84348
rect 65876 84346 65900 84348
rect 65956 84346 65962 84348
rect 65716 84294 65718 84346
rect 65898 84294 65900 84346
rect 65654 84292 65660 84294
rect 65716 84292 65740 84294
rect 65796 84292 65820 84294
rect 65876 84292 65900 84294
rect 65956 84292 65962 84294
rect 65654 84283 65962 84292
rect 96374 84348 96682 84357
rect 96374 84346 96380 84348
rect 96436 84346 96460 84348
rect 96516 84346 96540 84348
rect 96596 84346 96620 84348
rect 96676 84346 96682 84348
rect 96436 84294 96438 84346
rect 96618 84294 96620 84346
rect 96374 84292 96380 84294
rect 96436 84292 96460 84294
rect 96516 84292 96540 84294
rect 96596 84292 96620 84294
rect 96676 84292 96682 84294
rect 96374 84283 96682 84292
rect 66314 83804 66622 83813
rect 66314 83802 66320 83804
rect 66376 83802 66400 83804
rect 66456 83802 66480 83804
rect 66536 83802 66560 83804
rect 66616 83802 66622 83804
rect 66376 83750 66378 83802
rect 66558 83750 66560 83802
rect 66314 83748 66320 83750
rect 66376 83748 66400 83750
rect 66456 83748 66480 83750
rect 66536 83748 66560 83750
rect 66616 83748 66622 83750
rect 66314 83739 66622 83748
rect 97034 83804 97342 83813
rect 97034 83802 97040 83804
rect 97096 83802 97120 83804
rect 97176 83802 97200 83804
rect 97256 83802 97280 83804
rect 97336 83802 97342 83804
rect 97096 83750 97098 83802
rect 97278 83750 97280 83802
rect 97034 83748 97040 83750
rect 97096 83748 97120 83750
rect 97176 83748 97200 83750
rect 97256 83748 97280 83750
rect 97336 83748 97342 83750
rect 97034 83739 97342 83748
rect 65654 83260 65962 83269
rect 65654 83258 65660 83260
rect 65716 83258 65740 83260
rect 65796 83258 65820 83260
rect 65876 83258 65900 83260
rect 65956 83258 65962 83260
rect 65716 83206 65718 83258
rect 65898 83206 65900 83258
rect 65654 83204 65660 83206
rect 65716 83204 65740 83206
rect 65796 83204 65820 83206
rect 65876 83204 65900 83206
rect 65956 83204 65962 83206
rect 65654 83195 65962 83204
rect 96374 83260 96682 83269
rect 96374 83258 96380 83260
rect 96436 83258 96460 83260
rect 96516 83258 96540 83260
rect 96596 83258 96620 83260
rect 96676 83258 96682 83260
rect 96436 83206 96438 83258
rect 96618 83206 96620 83258
rect 96374 83204 96380 83206
rect 96436 83204 96460 83206
rect 96516 83204 96540 83206
rect 96596 83204 96620 83206
rect 96676 83204 96682 83206
rect 96374 83195 96682 83204
rect 66314 82716 66622 82725
rect 66314 82714 66320 82716
rect 66376 82714 66400 82716
rect 66456 82714 66480 82716
rect 66536 82714 66560 82716
rect 66616 82714 66622 82716
rect 66376 82662 66378 82714
rect 66558 82662 66560 82714
rect 66314 82660 66320 82662
rect 66376 82660 66400 82662
rect 66456 82660 66480 82662
rect 66536 82660 66560 82662
rect 66616 82660 66622 82662
rect 66314 82651 66622 82660
rect 97034 82716 97342 82725
rect 97034 82714 97040 82716
rect 97096 82714 97120 82716
rect 97176 82714 97200 82716
rect 97256 82714 97280 82716
rect 97336 82714 97342 82716
rect 97096 82662 97098 82714
rect 97278 82662 97280 82714
rect 97034 82660 97040 82662
rect 97096 82660 97120 82662
rect 97176 82660 97200 82662
rect 97256 82660 97280 82662
rect 97336 82660 97342 82662
rect 97034 82651 97342 82660
rect 65654 82172 65962 82181
rect 65654 82170 65660 82172
rect 65716 82170 65740 82172
rect 65796 82170 65820 82172
rect 65876 82170 65900 82172
rect 65956 82170 65962 82172
rect 65716 82118 65718 82170
rect 65898 82118 65900 82170
rect 65654 82116 65660 82118
rect 65716 82116 65740 82118
rect 65796 82116 65820 82118
rect 65876 82116 65900 82118
rect 65956 82116 65962 82118
rect 65654 82107 65962 82116
rect 96374 82172 96682 82181
rect 96374 82170 96380 82172
rect 96436 82170 96460 82172
rect 96516 82170 96540 82172
rect 96596 82170 96620 82172
rect 96676 82170 96682 82172
rect 96436 82118 96438 82170
rect 96618 82118 96620 82170
rect 96374 82116 96380 82118
rect 96436 82116 96460 82118
rect 96516 82116 96540 82118
rect 96596 82116 96620 82118
rect 96676 82116 96682 82118
rect 96374 82107 96682 82116
rect 66314 81628 66622 81637
rect 66314 81626 66320 81628
rect 66376 81626 66400 81628
rect 66456 81626 66480 81628
rect 66536 81626 66560 81628
rect 66616 81626 66622 81628
rect 66376 81574 66378 81626
rect 66558 81574 66560 81626
rect 66314 81572 66320 81574
rect 66376 81572 66400 81574
rect 66456 81572 66480 81574
rect 66536 81572 66560 81574
rect 66616 81572 66622 81574
rect 66314 81563 66622 81572
rect 97034 81628 97342 81637
rect 97034 81626 97040 81628
rect 97096 81626 97120 81628
rect 97176 81626 97200 81628
rect 97256 81626 97280 81628
rect 97336 81626 97342 81628
rect 97096 81574 97098 81626
rect 97278 81574 97280 81626
rect 97034 81572 97040 81574
rect 97096 81572 97120 81574
rect 97176 81572 97200 81574
rect 97256 81572 97280 81574
rect 97336 81572 97342 81574
rect 97034 81563 97342 81572
rect 65654 81084 65962 81093
rect 65654 81082 65660 81084
rect 65716 81082 65740 81084
rect 65796 81082 65820 81084
rect 65876 81082 65900 81084
rect 65956 81082 65962 81084
rect 65716 81030 65718 81082
rect 65898 81030 65900 81082
rect 65654 81028 65660 81030
rect 65716 81028 65740 81030
rect 65796 81028 65820 81030
rect 65876 81028 65900 81030
rect 65956 81028 65962 81030
rect 65654 81019 65962 81028
rect 96374 81084 96682 81093
rect 96374 81082 96380 81084
rect 96436 81082 96460 81084
rect 96516 81082 96540 81084
rect 96596 81082 96620 81084
rect 96676 81082 96682 81084
rect 96436 81030 96438 81082
rect 96618 81030 96620 81082
rect 96374 81028 96380 81030
rect 96436 81028 96460 81030
rect 96516 81028 96540 81030
rect 96596 81028 96620 81030
rect 96676 81028 96682 81030
rect 96374 81019 96682 81028
rect 66314 80540 66622 80549
rect 66314 80538 66320 80540
rect 66376 80538 66400 80540
rect 66456 80538 66480 80540
rect 66536 80538 66560 80540
rect 66616 80538 66622 80540
rect 66376 80486 66378 80538
rect 66558 80486 66560 80538
rect 66314 80484 66320 80486
rect 66376 80484 66400 80486
rect 66456 80484 66480 80486
rect 66536 80484 66560 80486
rect 66616 80484 66622 80486
rect 66314 80475 66622 80484
rect 97034 80540 97342 80549
rect 97034 80538 97040 80540
rect 97096 80538 97120 80540
rect 97176 80538 97200 80540
rect 97256 80538 97280 80540
rect 97336 80538 97342 80540
rect 97096 80486 97098 80538
rect 97278 80486 97280 80538
rect 97034 80484 97040 80486
rect 97096 80484 97120 80486
rect 97176 80484 97200 80486
rect 97256 80484 97280 80486
rect 97336 80484 97342 80486
rect 97034 80475 97342 80484
rect 65654 79996 65962 80005
rect 65654 79994 65660 79996
rect 65716 79994 65740 79996
rect 65796 79994 65820 79996
rect 65876 79994 65900 79996
rect 65956 79994 65962 79996
rect 65716 79942 65718 79994
rect 65898 79942 65900 79994
rect 65654 79940 65660 79942
rect 65716 79940 65740 79942
rect 65796 79940 65820 79942
rect 65876 79940 65900 79942
rect 65956 79940 65962 79942
rect 65654 79931 65962 79940
rect 96374 79996 96682 80005
rect 96374 79994 96380 79996
rect 96436 79994 96460 79996
rect 96516 79994 96540 79996
rect 96596 79994 96620 79996
rect 96676 79994 96682 79996
rect 96436 79942 96438 79994
rect 96618 79942 96620 79994
rect 96374 79940 96380 79942
rect 96436 79940 96460 79942
rect 96516 79940 96540 79942
rect 96596 79940 96620 79942
rect 96676 79940 96682 79942
rect 96374 79931 96682 79940
rect 66314 79452 66622 79461
rect 66314 79450 66320 79452
rect 66376 79450 66400 79452
rect 66456 79450 66480 79452
rect 66536 79450 66560 79452
rect 66616 79450 66622 79452
rect 66376 79398 66378 79450
rect 66558 79398 66560 79450
rect 66314 79396 66320 79398
rect 66376 79396 66400 79398
rect 66456 79396 66480 79398
rect 66536 79396 66560 79398
rect 66616 79396 66622 79398
rect 66314 79387 66622 79396
rect 97034 79452 97342 79461
rect 97034 79450 97040 79452
rect 97096 79450 97120 79452
rect 97176 79450 97200 79452
rect 97256 79450 97280 79452
rect 97336 79450 97342 79452
rect 97096 79398 97098 79450
rect 97278 79398 97280 79450
rect 97034 79396 97040 79398
rect 97096 79396 97120 79398
rect 97176 79396 97200 79398
rect 97256 79396 97280 79398
rect 97336 79396 97342 79398
rect 97034 79387 97342 79396
rect 65654 78908 65962 78917
rect 65654 78906 65660 78908
rect 65716 78906 65740 78908
rect 65796 78906 65820 78908
rect 65876 78906 65900 78908
rect 65956 78906 65962 78908
rect 65716 78854 65718 78906
rect 65898 78854 65900 78906
rect 65654 78852 65660 78854
rect 65716 78852 65740 78854
rect 65796 78852 65820 78854
rect 65876 78852 65900 78854
rect 65956 78852 65962 78854
rect 65654 78843 65962 78852
rect 96374 78908 96682 78917
rect 96374 78906 96380 78908
rect 96436 78906 96460 78908
rect 96516 78906 96540 78908
rect 96596 78906 96620 78908
rect 96676 78906 96682 78908
rect 96436 78854 96438 78906
rect 96618 78854 96620 78906
rect 96374 78852 96380 78854
rect 96436 78852 96460 78854
rect 96516 78852 96540 78854
rect 96596 78852 96620 78854
rect 96676 78852 96682 78854
rect 96374 78843 96682 78852
rect 66314 78364 66622 78373
rect 66314 78362 66320 78364
rect 66376 78362 66400 78364
rect 66456 78362 66480 78364
rect 66536 78362 66560 78364
rect 66616 78362 66622 78364
rect 66376 78310 66378 78362
rect 66558 78310 66560 78362
rect 66314 78308 66320 78310
rect 66376 78308 66400 78310
rect 66456 78308 66480 78310
rect 66536 78308 66560 78310
rect 66616 78308 66622 78310
rect 66314 78299 66622 78308
rect 97034 78364 97342 78373
rect 97034 78362 97040 78364
rect 97096 78362 97120 78364
rect 97176 78362 97200 78364
rect 97256 78362 97280 78364
rect 97336 78362 97342 78364
rect 97096 78310 97098 78362
rect 97278 78310 97280 78362
rect 97034 78308 97040 78310
rect 97096 78308 97120 78310
rect 97176 78308 97200 78310
rect 97256 78308 97280 78310
rect 97336 78308 97342 78310
rect 97034 78299 97342 78308
rect 65654 77820 65962 77829
rect 65654 77818 65660 77820
rect 65716 77818 65740 77820
rect 65796 77818 65820 77820
rect 65876 77818 65900 77820
rect 65956 77818 65962 77820
rect 65716 77766 65718 77818
rect 65898 77766 65900 77818
rect 65654 77764 65660 77766
rect 65716 77764 65740 77766
rect 65796 77764 65820 77766
rect 65876 77764 65900 77766
rect 65956 77764 65962 77766
rect 65654 77755 65962 77764
rect 96374 77820 96682 77829
rect 96374 77818 96380 77820
rect 96436 77818 96460 77820
rect 96516 77818 96540 77820
rect 96596 77818 96620 77820
rect 96676 77818 96682 77820
rect 96436 77766 96438 77818
rect 96618 77766 96620 77818
rect 96374 77764 96380 77766
rect 96436 77764 96460 77766
rect 96516 77764 96540 77766
rect 96596 77764 96620 77766
rect 96676 77764 96682 77766
rect 96374 77755 96682 77764
rect 53104 77716 53156 77722
rect 53104 77658 53156 77664
rect 55128 77716 55180 77722
rect 55128 77658 55180 77664
rect 57336 77716 57388 77722
rect 57336 77658 57388 77664
rect 59176 77716 59228 77722
rect 59176 77658 59228 77664
rect 51264 77444 51316 77450
rect 51264 77386 51316 77392
rect 53380 77444 53432 77450
rect 53380 77386 53432 77392
rect 55588 77444 55640 77450
rect 55588 77386 55640 77392
rect 57428 77444 57480 77450
rect 57428 77386 57480 77392
rect 59268 77444 59320 77450
rect 59268 77386 59320 77392
rect 51172 77172 51224 77178
rect 51172 77114 51224 77120
rect 51276 76838 51304 77386
rect 53288 77376 53340 77382
rect 53288 77318 53340 77324
rect 53196 77104 53248 77110
rect 53196 77046 53248 77052
rect 51264 76832 51316 76838
rect 51264 76774 51316 76780
rect 49976 74996 50028 75002
rect 49976 74938 50028 74944
rect 51080 74996 51132 75002
rect 51080 74938 51132 74944
rect 51276 71913 51304 76774
rect 53208 75002 53236 77046
rect 53300 76838 53328 77318
rect 53288 76832 53340 76838
rect 53288 76774 53340 76780
rect 53300 75857 53328 76774
rect 53286 75848 53342 75857
rect 53286 75783 53342 75792
rect 53392 75002 53420 77386
rect 55600 76838 55628 77386
rect 56876 77376 56928 77382
rect 56876 77318 56928 77324
rect 55588 76832 55640 76838
rect 55588 76774 55640 76780
rect 53196 74996 53248 75002
rect 53196 74938 53248 74944
rect 53380 74996 53432 75002
rect 53380 74938 53432 74944
rect 55600 74633 55628 76774
rect 56888 75002 56916 77318
rect 57440 75002 57468 77386
rect 57520 77376 57572 77382
rect 57520 77318 57572 77324
rect 57532 76838 57560 77318
rect 57520 76832 57572 76838
rect 57520 76774 57572 76780
rect 56876 74996 56928 75002
rect 56876 74938 56928 74944
rect 57428 74996 57480 75002
rect 57428 74938 57480 74944
rect 55586 74624 55642 74633
rect 55586 74559 55642 74568
rect 57532 73953 57560 76774
rect 59280 75002 59308 77386
rect 66314 77276 66622 77285
rect 66314 77274 66320 77276
rect 66376 77274 66400 77276
rect 66456 77274 66480 77276
rect 66536 77274 66560 77276
rect 66616 77274 66622 77276
rect 66376 77222 66378 77274
rect 66558 77222 66560 77274
rect 66314 77220 66320 77222
rect 66376 77220 66400 77222
rect 66456 77220 66480 77222
rect 66536 77220 66560 77222
rect 66616 77220 66622 77222
rect 66314 77211 66622 77220
rect 97034 77276 97342 77285
rect 97034 77274 97040 77276
rect 97096 77274 97120 77276
rect 97176 77274 97200 77276
rect 97256 77274 97280 77276
rect 97336 77274 97342 77276
rect 97096 77222 97098 77274
rect 97278 77222 97280 77274
rect 97034 77220 97040 77222
rect 97096 77220 97120 77222
rect 97176 77220 97200 77222
rect 97256 77220 97280 77222
rect 97336 77220 97342 77222
rect 97034 77211 97342 77220
rect 65654 76732 65962 76741
rect 65654 76730 65660 76732
rect 65716 76730 65740 76732
rect 65796 76730 65820 76732
rect 65876 76730 65900 76732
rect 65956 76730 65962 76732
rect 65716 76678 65718 76730
rect 65898 76678 65900 76730
rect 65654 76676 65660 76678
rect 65716 76676 65740 76678
rect 65796 76676 65820 76678
rect 65876 76676 65900 76678
rect 65956 76676 65962 76678
rect 65654 76667 65962 76676
rect 96374 76732 96682 76741
rect 96374 76730 96380 76732
rect 96436 76730 96460 76732
rect 96516 76730 96540 76732
rect 96596 76730 96620 76732
rect 96676 76730 96682 76732
rect 96436 76678 96438 76730
rect 96618 76678 96620 76730
rect 96374 76676 96380 76678
rect 96436 76676 96460 76678
rect 96516 76676 96540 76678
rect 96596 76676 96620 76678
rect 96676 76676 96682 76678
rect 96374 76667 96682 76676
rect 66314 76188 66622 76197
rect 66314 76186 66320 76188
rect 66376 76186 66400 76188
rect 66456 76186 66480 76188
rect 66536 76186 66560 76188
rect 66616 76186 66622 76188
rect 66376 76134 66378 76186
rect 66558 76134 66560 76186
rect 66314 76132 66320 76134
rect 66376 76132 66400 76134
rect 66456 76132 66480 76134
rect 66536 76132 66560 76134
rect 66616 76132 66622 76134
rect 66314 76123 66622 76132
rect 97034 76188 97342 76197
rect 97034 76186 97040 76188
rect 97096 76186 97120 76188
rect 97176 76186 97200 76188
rect 97256 76186 97280 76188
rect 97336 76186 97342 76188
rect 97096 76134 97098 76186
rect 97278 76134 97280 76186
rect 97034 76132 97040 76134
rect 97096 76132 97120 76134
rect 97176 76132 97200 76134
rect 97256 76132 97280 76134
rect 97336 76132 97342 76134
rect 97034 76123 97342 76132
rect 65654 75644 65962 75653
rect 65654 75642 65660 75644
rect 65716 75642 65740 75644
rect 65796 75642 65820 75644
rect 65876 75642 65900 75644
rect 65956 75642 65962 75644
rect 65716 75590 65718 75642
rect 65898 75590 65900 75642
rect 65654 75588 65660 75590
rect 65716 75588 65740 75590
rect 65796 75588 65820 75590
rect 65876 75588 65900 75590
rect 65956 75588 65962 75590
rect 65654 75579 65962 75588
rect 96374 75644 96682 75653
rect 96374 75642 96380 75644
rect 96436 75642 96460 75644
rect 96516 75642 96540 75644
rect 96596 75642 96620 75644
rect 96676 75642 96682 75644
rect 96436 75590 96438 75642
rect 96618 75590 96620 75642
rect 96374 75588 96380 75590
rect 96436 75588 96460 75590
rect 96516 75588 96540 75590
rect 96596 75588 96620 75590
rect 96676 75588 96682 75590
rect 96374 75579 96682 75588
rect 66314 75100 66622 75109
rect 66314 75098 66320 75100
rect 66376 75098 66400 75100
rect 66456 75098 66480 75100
rect 66536 75098 66560 75100
rect 66616 75098 66622 75100
rect 66376 75046 66378 75098
rect 66558 75046 66560 75098
rect 66314 75044 66320 75046
rect 66376 75044 66400 75046
rect 66456 75044 66480 75046
rect 66536 75044 66560 75046
rect 66616 75044 66622 75046
rect 66314 75035 66622 75044
rect 97034 75100 97342 75109
rect 97034 75098 97040 75100
rect 97096 75098 97120 75100
rect 97176 75098 97200 75100
rect 97256 75098 97280 75100
rect 97336 75098 97342 75100
rect 97096 75046 97098 75098
rect 97278 75046 97280 75098
rect 97034 75044 97040 75046
rect 97096 75044 97120 75046
rect 97176 75044 97200 75046
rect 97256 75044 97280 75046
rect 97336 75044 97342 75046
rect 97034 75035 97342 75044
rect 59268 74996 59320 75002
rect 59268 74938 59320 74944
rect 83924 74860 83976 74866
rect 83924 74802 83976 74808
rect 65654 74556 65962 74565
rect 65654 74554 65660 74556
rect 65716 74554 65740 74556
rect 65796 74554 65820 74556
rect 65876 74554 65900 74556
rect 65956 74554 65962 74556
rect 65716 74502 65718 74554
rect 65898 74502 65900 74554
rect 65654 74500 65660 74502
rect 65716 74500 65740 74502
rect 65796 74500 65820 74502
rect 65876 74500 65900 74502
rect 65956 74500 65962 74502
rect 65654 74491 65962 74500
rect 66314 74012 66622 74021
rect 66314 74010 66320 74012
rect 66376 74010 66400 74012
rect 66456 74010 66480 74012
rect 66536 74010 66560 74012
rect 66616 74010 66622 74012
rect 66376 73958 66378 74010
rect 66558 73958 66560 74010
rect 66314 73956 66320 73958
rect 66376 73956 66400 73958
rect 66456 73956 66480 73958
rect 66536 73956 66560 73958
rect 66616 73956 66622 73958
rect 57518 73944 57574 73953
rect 66314 73947 66622 73956
rect 57518 73879 57574 73888
rect 65654 73468 65962 73477
rect 65654 73466 65660 73468
rect 65716 73466 65740 73468
rect 65796 73466 65820 73468
rect 65876 73466 65900 73468
rect 65956 73466 65962 73468
rect 65716 73414 65718 73466
rect 65898 73414 65900 73466
rect 65654 73412 65660 73414
rect 65716 73412 65740 73414
rect 65796 73412 65820 73414
rect 65876 73412 65900 73414
rect 65956 73412 65962 73414
rect 65654 73403 65962 73412
rect 66314 72924 66622 72933
rect 66314 72922 66320 72924
rect 66376 72922 66400 72924
rect 66456 72922 66480 72924
rect 66536 72922 66560 72924
rect 66616 72922 66622 72924
rect 66376 72870 66378 72922
rect 66558 72870 66560 72922
rect 66314 72868 66320 72870
rect 66376 72868 66400 72870
rect 66456 72868 66480 72870
rect 66536 72868 66560 72870
rect 66616 72868 66622 72870
rect 66314 72859 66622 72868
rect 65654 72380 65962 72389
rect 65654 72378 65660 72380
rect 65716 72378 65740 72380
rect 65796 72378 65820 72380
rect 65876 72378 65900 72380
rect 65956 72378 65962 72380
rect 65716 72326 65718 72378
rect 65898 72326 65900 72378
rect 65654 72324 65660 72326
rect 65716 72324 65740 72326
rect 65796 72324 65820 72326
rect 65876 72324 65900 72326
rect 65956 72324 65962 72326
rect 65654 72315 65962 72324
rect 51262 71904 51318 71913
rect 51262 71839 51318 71848
rect 66314 71836 66622 71845
rect 66314 71834 66320 71836
rect 66376 71834 66400 71836
rect 66456 71834 66480 71836
rect 66536 71834 66560 71836
rect 66616 71834 66622 71836
rect 66376 71782 66378 71834
rect 66558 71782 66560 71834
rect 66314 71780 66320 71782
rect 66376 71780 66400 71782
rect 66456 71780 66480 71782
rect 66536 71780 66560 71782
rect 66616 71780 66622 71782
rect 66314 71771 66622 71780
rect 65654 71292 65962 71301
rect 65654 71290 65660 71292
rect 65716 71290 65740 71292
rect 65796 71290 65820 71292
rect 65876 71290 65900 71292
rect 65956 71290 65962 71292
rect 65716 71238 65718 71290
rect 65898 71238 65900 71290
rect 65654 71236 65660 71238
rect 65716 71236 65740 71238
rect 65796 71236 65820 71238
rect 65876 71236 65900 71238
rect 65956 71236 65962 71238
rect 65654 71227 65962 71236
rect 66314 70748 66622 70757
rect 66314 70746 66320 70748
rect 66376 70746 66400 70748
rect 66456 70746 66480 70748
rect 66536 70746 66560 70748
rect 66616 70746 66622 70748
rect 66376 70694 66378 70746
rect 66558 70694 66560 70746
rect 66314 70692 66320 70694
rect 66376 70692 66400 70694
rect 66456 70692 66480 70694
rect 66536 70692 66560 70694
rect 66616 70692 66622 70694
rect 66314 70683 66622 70692
rect 65654 70204 65962 70213
rect 65654 70202 65660 70204
rect 65716 70202 65740 70204
rect 65796 70202 65820 70204
rect 65876 70202 65900 70204
rect 65956 70202 65962 70204
rect 65716 70150 65718 70202
rect 65898 70150 65900 70202
rect 65654 70148 65660 70150
rect 65716 70148 65740 70150
rect 65796 70148 65820 70150
rect 65876 70148 65900 70150
rect 65956 70148 65962 70150
rect 65654 70139 65962 70148
rect 66314 69660 66622 69669
rect 66314 69658 66320 69660
rect 66376 69658 66400 69660
rect 66456 69658 66480 69660
rect 66536 69658 66560 69660
rect 66616 69658 66622 69660
rect 66376 69606 66378 69658
rect 66558 69606 66560 69658
rect 66314 69604 66320 69606
rect 66376 69604 66400 69606
rect 66456 69604 66480 69606
rect 66536 69604 66560 69606
rect 66616 69604 66622 69606
rect 66314 69595 66622 69604
rect 65654 69116 65962 69125
rect 65654 69114 65660 69116
rect 65716 69114 65740 69116
rect 65796 69114 65820 69116
rect 65876 69114 65900 69116
rect 65956 69114 65962 69116
rect 65716 69062 65718 69114
rect 65898 69062 65900 69114
rect 65654 69060 65660 69062
rect 65716 69060 65740 69062
rect 65796 69060 65820 69062
rect 65876 69060 65900 69062
rect 65956 69060 65962 69062
rect 65654 69051 65962 69060
rect 66314 68572 66622 68581
rect 66314 68570 66320 68572
rect 66376 68570 66400 68572
rect 66456 68570 66480 68572
rect 66536 68570 66560 68572
rect 66616 68570 66622 68572
rect 66376 68518 66378 68570
rect 66558 68518 66560 68570
rect 66314 68516 66320 68518
rect 66376 68516 66400 68518
rect 66456 68516 66480 68518
rect 66536 68516 66560 68518
rect 66616 68516 66622 68518
rect 66314 68507 66622 68516
rect 65654 68028 65962 68037
rect 65654 68026 65660 68028
rect 65716 68026 65740 68028
rect 65796 68026 65820 68028
rect 65876 68026 65900 68028
rect 65956 68026 65962 68028
rect 65716 67974 65718 68026
rect 65898 67974 65900 68026
rect 65654 67972 65660 67974
rect 65716 67972 65740 67974
rect 65796 67972 65820 67974
rect 65876 67972 65900 67974
rect 65956 67972 65962 67974
rect 65654 67963 65962 67972
rect 66314 67484 66622 67493
rect 66314 67482 66320 67484
rect 66376 67482 66400 67484
rect 66456 67482 66480 67484
rect 66536 67482 66560 67484
rect 66616 67482 66622 67484
rect 66376 67430 66378 67482
rect 66558 67430 66560 67482
rect 66314 67428 66320 67430
rect 66376 67428 66400 67430
rect 66456 67428 66480 67430
rect 66536 67428 66560 67430
rect 66616 67428 66622 67430
rect 66314 67419 66622 67428
rect 65654 66940 65962 66949
rect 65654 66938 65660 66940
rect 65716 66938 65740 66940
rect 65796 66938 65820 66940
rect 65876 66938 65900 66940
rect 65956 66938 65962 66940
rect 65716 66886 65718 66938
rect 65898 66886 65900 66938
rect 65654 66884 65660 66886
rect 65716 66884 65740 66886
rect 65796 66884 65820 66886
rect 65876 66884 65900 66886
rect 65956 66884 65962 66886
rect 65654 66875 65962 66884
rect 66314 66396 66622 66405
rect 66314 66394 66320 66396
rect 66376 66394 66400 66396
rect 66456 66394 66480 66396
rect 66536 66394 66560 66396
rect 66616 66394 66622 66396
rect 66376 66342 66378 66394
rect 66558 66342 66560 66394
rect 66314 66340 66320 66342
rect 66376 66340 66400 66342
rect 66456 66340 66480 66342
rect 66536 66340 66560 66342
rect 66616 66340 66622 66342
rect 66314 66331 66622 66340
rect 65654 65852 65962 65861
rect 65654 65850 65660 65852
rect 65716 65850 65740 65852
rect 65796 65850 65820 65852
rect 65876 65850 65900 65852
rect 65956 65850 65962 65852
rect 65716 65798 65718 65850
rect 65898 65798 65900 65850
rect 65654 65796 65660 65798
rect 65716 65796 65740 65798
rect 65796 65796 65820 65798
rect 65876 65796 65900 65798
rect 65956 65796 65962 65798
rect 65654 65787 65962 65796
rect 66314 65308 66622 65317
rect 66314 65306 66320 65308
rect 66376 65306 66400 65308
rect 66456 65306 66480 65308
rect 66536 65306 66560 65308
rect 66616 65306 66622 65308
rect 66376 65254 66378 65306
rect 66558 65254 66560 65306
rect 66314 65252 66320 65254
rect 66376 65252 66400 65254
rect 66456 65252 66480 65254
rect 66536 65252 66560 65254
rect 66616 65252 66622 65254
rect 66314 65243 66622 65252
rect 65654 64764 65962 64773
rect 65654 64762 65660 64764
rect 65716 64762 65740 64764
rect 65796 64762 65820 64764
rect 65876 64762 65900 64764
rect 65956 64762 65962 64764
rect 65716 64710 65718 64762
rect 65898 64710 65900 64762
rect 65654 64708 65660 64710
rect 65716 64708 65740 64710
rect 65796 64708 65820 64710
rect 65876 64708 65900 64710
rect 65956 64708 65962 64710
rect 65654 64699 65962 64708
rect 66314 64220 66622 64229
rect 66314 64218 66320 64220
rect 66376 64218 66400 64220
rect 66456 64218 66480 64220
rect 66536 64218 66560 64220
rect 66616 64218 66622 64220
rect 66376 64166 66378 64218
rect 66558 64166 66560 64218
rect 66314 64164 66320 64166
rect 66376 64164 66400 64166
rect 66456 64164 66480 64166
rect 66536 64164 66560 64166
rect 66616 64164 66622 64166
rect 66314 64155 66622 64164
rect 65654 63676 65962 63685
rect 65654 63674 65660 63676
rect 65716 63674 65740 63676
rect 65796 63674 65820 63676
rect 65876 63674 65900 63676
rect 65956 63674 65962 63676
rect 65716 63622 65718 63674
rect 65898 63622 65900 63674
rect 65654 63620 65660 63622
rect 65716 63620 65740 63622
rect 65796 63620 65820 63622
rect 65876 63620 65900 63622
rect 65956 63620 65962 63622
rect 65654 63611 65962 63620
rect 66314 63132 66622 63141
rect 66314 63130 66320 63132
rect 66376 63130 66400 63132
rect 66456 63130 66480 63132
rect 66536 63130 66560 63132
rect 66616 63130 66622 63132
rect 66376 63078 66378 63130
rect 66558 63078 66560 63130
rect 66314 63076 66320 63078
rect 66376 63076 66400 63078
rect 66456 63076 66480 63078
rect 66536 63076 66560 63078
rect 66616 63076 66622 63078
rect 66314 63067 66622 63076
rect 65654 62588 65962 62597
rect 65654 62586 65660 62588
rect 65716 62586 65740 62588
rect 65796 62586 65820 62588
rect 65876 62586 65900 62588
rect 65956 62586 65962 62588
rect 65716 62534 65718 62586
rect 65898 62534 65900 62586
rect 65654 62532 65660 62534
rect 65716 62532 65740 62534
rect 65796 62532 65820 62534
rect 65876 62532 65900 62534
rect 65956 62532 65962 62534
rect 65654 62523 65962 62532
rect 66314 62044 66622 62053
rect 66314 62042 66320 62044
rect 66376 62042 66400 62044
rect 66456 62042 66480 62044
rect 66536 62042 66560 62044
rect 66616 62042 66622 62044
rect 66376 61990 66378 62042
rect 66558 61990 66560 62042
rect 66314 61988 66320 61990
rect 66376 61988 66400 61990
rect 66456 61988 66480 61990
rect 66536 61988 66560 61990
rect 66616 61988 66622 61990
rect 66314 61979 66622 61988
rect 65654 61500 65962 61509
rect 65654 61498 65660 61500
rect 65716 61498 65740 61500
rect 65796 61498 65820 61500
rect 65876 61498 65900 61500
rect 65956 61498 65962 61500
rect 65716 61446 65718 61498
rect 65898 61446 65900 61498
rect 65654 61444 65660 61446
rect 65716 61444 65740 61446
rect 65796 61444 65820 61446
rect 65876 61444 65900 61446
rect 65956 61444 65962 61446
rect 65654 61435 65962 61444
rect 77116 61396 77168 61402
rect 77116 61338 77168 61344
rect 82452 61396 82504 61402
rect 82452 61338 82504 61344
rect 77024 61192 77076 61198
rect 77024 61134 77076 61140
rect 71780 61056 71832 61062
rect 71780 60998 71832 61004
rect 66314 60956 66622 60965
rect 66314 60954 66320 60956
rect 66376 60954 66400 60956
rect 66456 60954 66480 60956
rect 66536 60954 66560 60956
rect 66616 60954 66622 60956
rect 66376 60902 66378 60954
rect 66558 60902 66560 60954
rect 66314 60900 66320 60902
rect 66376 60900 66400 60902
rect 66456 60900 66480 60902
rect 66536 60900 66560 60902
rect 66616 60900 66622 60902
rect 66314 60891 66622 60900
rect 48412 60784 48464 60790
rect 48412 60726 48464 60732
rect 49424 60784 49476 60790
rect 49424 60726 49476 60732
rect 28816 60716 28868 60722
rect 28816 60658 28868 60664
rect 46664 60716 46716 60722
rect 46664 60658 46716 60664
rect 34934 60412 35242 60421
rect 34934 60410 34940 60412
rect 34996 60410 35020 60412
rect 35076 60410 35100 60412
rect 35156 60410 35180 60412
rect 35236 60410 35242 60412
rect 34996 60358 34998 60410
rect 35178 60358 35180 60410
rect 34934 60356 34940 60358
rect 34996 60356 35020 60358
rect 35076 60356 35100 60358
rect 35156 60356 35180 60358
rect 35236 60356 35242 60358
rect 34934 60347 35242 60356
rect 48424 60314 48452 60726
rect 65654 60412 65962 60421
rect 65654 60410 65660 60412
rect 65716 60410 65740 60412
rect 65796 60410 65820 60412
rect 65876 60410 65900 60412
rect 65956 60410 65962 60412
rect 65716 60358 65718 60410
rect 65898 60358 65900 60410
rect 65654 60356 65660 60358
rect 65716 60356 65740 60358
rect 65796 60356 65820 60358
rect 65876 60356 65900 60358
rect 65956 60356 65962 60358
rect 65654 60347 65962 60356
rect 29184 60308 29236 60314
rect 29184 60250 29236 60256
rect 48412 60308 48464 60314
rect 48412 60250 48464 60256
rect 29196 58177 29224 60250
rect 57060 60036 57112 60042
rect 57060 59978 57112 59984
rect 35594 59868 35902 59877
rect 35594 59866 35600 59868
rect 35656 59866 35680 59868
rect 35736 59866 35760 59868
rect 35816 59866 35840 59868
rect 35896 59866 35902 59868
rect 35656 59814 35658 59866
rect 35838 59814 35840 59866
rect 35594 59812 35600 59814
rect 35656 59812 35680 59814
rect 35736 59812 35760 59814
rect 35816 59812 35840 59814
rect 35896 59812 35902 59814
rect 35594 59803 35902 59812
rect 57072 58682 57100 59978
rect 66314 59868 66622 59877
rect 66314 59866 66320 59868
rect 66376 59866 66400 59868
rect 66456 59866 66480 59868
rect 66536 59866 66560 59868
rect 66616 59866 66622 59868
rect 66376 59814 66378 59866
rect 66558 59814 66560 59866
rect 66314 59812 66320 59814
rect 66376 59812 66400 59814
rect 66456 59812 66480 59814
rect 66536 59812 66560 59814
rect 66616 59812 66622 59814
rect 66314 59803 66622 59812
rect 71792 58857 71820 60998
rect 77036 60178 77064 61134
rect 77128 60761 77156 61338
rect 79692 61260 79744 61266
rect 79692 61202 79744 61208
rect 79876 61260 79928 61266
rect 79876 61202 79928 61208
rect 77760 61124 77812 61130
rect 77760 61066 77812 61072
rect 79140 61124 79192 61130
rect 79140 61066 79192 61072
rect 79600 61124 79652 61130
rect 79600 61066 79652 61072
rect 77114 60752 77170 60761
rect 77114 60687 77170 60696
rect 77772 60654 77800 61066
rect 79152 60858 79180 61066
rect 79140 60852 79192 60858
rect 79140 60794 79192 60800
rect 77760 60648 77812 60654
rect 77760 60590 77812 60596
rect 77024 60172 77076 60178
rect 77024 60114 77076 60120
rect 71778 58848 71834 58857
rect 71778 58783 71834 58792
rect 57060 58676 57112 58682
rect 57060 58618 57112 58624
rect 79152 58585 79180 60794
rect 79232 60716 79284 60722
rect 79232 60658 79284 60664
rect 79244 60110 79272 60658
rect 79612 60654 79640 61066
rect 79704 60722 79732 61202
rect 79888 60858 79916 61202
rect 81532 61192 81584 61198
rect 81532 61134 81584 61140
rect 79876 60852 79928 60858
rect 79876 60794 79928 60800
rect 79692 60716 79744 60722
rect 79692 60658 79744 60664
rect 79600 60648 79652 60654
rect 79600 60590 79652 60596
rect 79704 60518 79732 60658
rect 81544 60654 81572 61134
rect 82464 61130 82492 61338
rect 83936 61198 83964 74802
rect 96374 74556 96682 74565
rect 96374 74554 96380 74556
rect 96436 74554 96460 74556
rect 96516 74554 96540 74556
rect 96596 74554 96620 74556
rect 96676 74554 96682 74556
rect 96436 74502 96438 74554
rect 96618 74502 96620 74554
rect 96374 74500 96380 74502
rect 96436 74500 96460 74502
rect 96516 74500 96540 74502
rect 96596 74500 96620 74502
rect 96676 74500 96682 74502
rect 96374 74491 96682 74500
rect 97034 74012 97342 74021
rect 97034 74010 97040 74012
rect 97096 74010 97120 74012
rect 97176 74010 97200 74012
rect 97256 74010 97280 74012
rect 97336 74010 97342 74012
rect 97096 73958 97098 74010
rect 97278 73958 97280 74010
rect 97034 73956 97040 73958
rect 97096 73956 97120 73958
rect 97176 73956 97200 73958
rect 97256 73956 97280 73958
rect 97336 73956 97342 73958
rect 97034 73947 97342 73956
rect 96374 73468 96682 73477
rect 96374 73466 96380 73468
rect 96436 73466 96460 73468
rect 96516 73466 96540 73468
rect 96596 73466 96620 73468
rect 96676 73466 96682 73468
rect 96436 73414 96438 73466
rect 96618 73414 96620 73466
rect 96374 73412 96380 73414
rect 96436 73412 96460 73414
rect 96516 73412 96540 73414
rect 96596 73412 96620 73414
rect 96676 73412 96682 73414
rect 96374 73403 96682 73412
rect 97034 72924 97342 72933
rect 97034 72922 97040 72924
rect 97096 72922 97120 72924
rect 97176 72922 97200 72924
rect 97256 72922 97280 72924
rect 97336 72922 97342 72924
rect 97096 72870 97098 72922
rect 97278 72870 97280 72922
rect 97034 72868 97040 72870
rect 97096 72868 97120 72870
rect 97176 72868 97200 72870
rect 97256 72868 97280 72870
rect 97336 72868 97342 72870
rect 97034 72859 97342 72868
rect 96374 72380 96682 72389
rect 96374 72378 96380 72380
rect 96436 72378 96460 72380
rect 96516 72378 96540 72380
rect 96596 72378 96620 72380
rect 96676 72378 96682 72380
rect 96436 72326 96438 72378
rect 96618 72326 96620 72378
rect 96374 72324 96380 72326
rect 96436 72324 96460 72326
rect 96516 72324 96540 72326
rect 96596 72324 96620 72326
rect 96676 72324 96682 72326
rect 96374 72315 96682 72324
rect 97034 71836 97342 71845
rect 97034 71834 97040 71836
rect 97096 71834 97120 71836
rect 97176 71834 97200 71836
rect 97256 71834 97280 71836
rect 97336 71834 97342 71836
rect 97096 71782 97098 71834
rect 97278 71782 97280 71834
rect 97034 71780 97040 71782
rect 97096 71780 97120 71782
rect 97176 71780 97200 71782
rect 97256 71780 97280 71782
rect 97336 71780 97342 71782
rect 97034 71771 97342 71780
rect 96374 71292 96682 71301
rect 96374 71290 96380 71292
rect 96436 71290 96460 71292
rect 96516 71290 96540 71292
rect 96596 71290 96620 71292
rect 96676 71290 96682 71292
rect 96436 71238 96438 71290
rect 96618 71238 96620 71290
rect 96374 71236 96380 71238
rect 96436 71236 96460 71238
rect 96516 71236 96540 71238
rect 96596 71236 96620 71238
rect 96676 71236 96682 71238
rect 96374 71227 96682 71236
rect 97034 70748 97342 70757
rect 97034 70746 97040 70748
rect 97096 70746 97120 70748
rect 97176 70746 97200 70748
rect 97256 70746 97280 70748
rect 97336 70746 97342 70748
rect 97096 70694 97098 70746
rect 97278 70694 97280 70746
rect 97034 70692 97040 70694
rect 97096 70692 97120 70694
rect 97176 70692 97200 70694
rect 97256 70692 97280 70694
rect 97336 70692 97342 70694
rect 97034 70683 97342 70692
rect 96374 70204 96682 70213
rect 96374 70202 96380 70204
rect 96436 70202 96460 70204
rect 96516 70202 96540 70204
rect 96596 70202 96620 70204
rect 96676 70202 96682 70204
rect 96436 70150 96438 70202
rect 96618 70150 96620 70202
rect 96374 70148 96380 70150
rect 96436 70148 96460 70150
rect 96516 70148 96540 70150
rect 96596 70148 96620 70150
rect 96676 70148 96682 70150
rect 96374 70139 96682 70148
rect 97034 69660 97342 69669
rect 97034 69658 97040 69660
rect 97096 69658 97120 69660
rect 97176 69658 97200 69660
rect 97256 69658 97280 69660
rect 97336 69658 97342 69660
rect 97096 69606 97098 69658
rect 97278 69606 97280 69658
rect 97034 69604 97040 69606
rect 97096 69604 97120 69606
rect 97176 69604 97200 69606
rect 97256 69604 97280 69606
rect 97336 69604 97342 69606
rect 97034 69595 97342 69604
rect 96374 69116 96682 69125
rect 96374 69114 96380 69116
rect 96436 69114 96460 69116
rect 96516 69114 96540 69116
rect 96596 69114 96620 69116
rect 96676 69114 96682 69116
rect 96436 69062 96438 69114
rect 96618 69062 96620 69114
rect 96374 69060 96380 69062
rect 96436 69060 96460 69062
rect 96516 69060 96540 69062
rect 96596 69060 96620 69062
rect 96676 69060 96682 69062
rect 96374 69051 96682 69060
rect 97034 68572 97342 68581
rect 97034 68570 97040 68572
rect 97096 68570 97120 68572
rect 97176 68570 97200 68572
rect 97256 68570 97280 68572
rect 97336 68570 97342 68572
rect 97096 68518 97098 68570
rect 97278 68518 97280 68570
rect 97034 68516 97040 68518
rect 97096 68516 97120 68518
rect 97176 68516 97200 68518
rect 97256 68516 97280 68518
rect 97336 68516 97342 68518
rect 97034 68507 97342 68516
rect 96374 68028 96682 68037
rect 96374 68026 96380 68028
rect 96436 68026 96460 68028
rect 96516 68026 96540 68028
rect 96596 68026 96620 68028
rect 96676 68026 96682 68028
rect 96436 67974 96438 68026
rect 96618 67974 96620 68026
rect 96374 67972 96380 67974
rect 96436 67972 96460 67974
rect 96516 67972 96540 67974
rect 96596 67972 96620 67974
rect 96676 67972 96682 67974
rect 96374 67963 96682 67972
rect 97034 67484 97342 67493
rect 97034 67482 97040 67484
rect 97096 67482 97120 67484
rect 97176 67482 97200 67484
rect 97256 67482 97280 67484
rect 97336 67482 97342 67484
rect 97096 67430 97098 67482
rect 97278 67430 97280 67482
rect 97034 67428 97040 67430
rect 97096 67428 97120 67430
rect 97176 67428 97200 67430
rect 97256 67428 97280 67430
rect 97336 67428 97342 67430
rect 97034 67419 97342 67428
rect 96374 66940 96682 66949
rect 96374 66938 96380 66940
rect 96436 66938 96460 66940
rect 96516 66938 96540 66940
rect 96596 66938 96620 66940
rect 96676 66938 96682 66940
rect 96436 66886 96438 66938
rect 96618 66886 96620 66938
rect 96374 66884 96380 66886
rect 96436 66884 96460 66886
rect 96516 66884 96540 66886
rect 96596 66884 96620 66886
rect 96676 66884 96682 66886
rect 96374 66875 96682 66884
rect 97034 66396 97342 66405
rect 97034 66394 97040 66396
rect 97096 66394 97120 66396
rect 97176 66394 97200 66396
rect 97256 66394 97280 66396
rect 97336 66394 97342 66396
rect 97096 66342 97098 66394
rect 97278 66342 97280 66394
rect 97034 66340 97040 66342
rect 97096 66340 97120 66342
rect 97176 66340 97200 66342
rect 97256 66340 97280 66342
rect 97336 66340 97342 66342
rect 97034 66331 97342 66340
rect 96374 65852 96682 65861
rect 96374 65850 96380 65852
rect 96436 65850 96460 65852
rect 96516 65850 96540 65852
rect 96596 65850 96620 65852
rect 96676 65850 96682 65852
rect 96436 65798 96438 65850
rect 96618 65798 96620 65850
rect 96374 65796 96380 65798
rect 96436 65796 96460 65798
rect 96516 65796 96540 65798
rect 96596 65796 96620 65798
rect 96676 65796 96682 65798
rect 96374 65787 96682 65796
rect 97034 65308 97342 65317
rect 97034 65306 97040 65308
rect 97096 65306 97120 65308
rect 97176 65306 97200 65308
rect 97256 65306 97280 65308
rect 97336 65306 97342 65308
rect 97096 65254 97098 65306
rect 97278 65254 97280 65306
rect 97034 65252 97040 65254
rect 97096 65252 97120 65254
rect 97176 65252 97200 65254
rect 97256 65252 97280 65254
rect 97336 65252 97342 65254
rect 97034 65243 97342 65252
rect 96374 64764 96682 64773
rect 96374 64762 96380 64764
rect 96436 64762 96460 64764
rect 96516 64762 96540 64764
rect 96596 64762 96620 64764
rect 96676 64762 96682 64764
rect 96436 64710 96438 64762
rect 96618 64710 96620 64762
rect 96374 64708 96380 64710
rect 96436 64708 96460 64710
rect 96516 64708 96540 64710
rect 96596 64708 96620 64710
rect 96676 64708 96682 64710
rect 96374 64699 96682 64708
rect 97034 64220 97342 64229
rect 97034 64218 97040 64220
rect 97096 64218 97120 64220
rect 97176 64218 97200 64220
rect 97256 64218 97280 64220
rect 97336 64218 97342 64220
rect 97096 64166 97098 64218
rect 97278 64166 97280 64218
rect 97034 64164 97040 64166
rect 97096 64164 97120 64166
rect 97176 64164 97200 64166
rect 97256 64164 97280 64166
rect 97336 64164 97342 64166
rect 97034 64155 97342 64164
rect 96374 63676 96682 63685
rect 96374 63674 96380 63676
rect 96436 63674 96460 63676
rect 96516 63674 96540 63676
rect 96596 63674 96620 63676
rect 96676 63674 96682 63676
rect 96436 63622 96438 63674
rect 96618 63622 96620 63674
rect 96374 63620 96380 63622
rect 96436 63620 96460 63622
rect 96516 63620 96540 63622
rect 96596 63620 96620 63622
rect 96676 63620 96682 63622
rect 96374 63611 96682 63620
rect 97034 63132 97342 63141
rect 97034 63130 97040 63132
rect 97096 63130 97120 63132
rect 97176 63130 97200 63132
rect 97256 63130 97280 63132
rect 97336 63130 97342 63132
rect 97096 63078 97098 63130
rect 97278 63078 97280 63130
rect 97034 63076 97040 63078
rect 97096 63076 97120 63078
rect 97176 63076 97200 63078
rect 97256 63076 97280 63078
rect 97336 63076 97342 63078
rect 97034 63067 97342 63076
rect 96252 62892 96304 62898
rect 96252 62834 96304 62840
rect 96264 61402 96292 62834
rect 100392 62688 100444 62694
rect 100390 62656 100392 62665
rect 100444 62656 100446 62665
rect 96374 62588 96682 62597
rect 100390 62591 100446 62600
rect 96374 62586 96380 62588
rect 96436 62586 96460 62588
rect 96516 62586 96540 62588
rect 96596 62586 96620 62588
rect 96676 62586 96682 62588
rect 96436 62534 96438 62586
rect 96618 62534 96620 62586
rect 96374 62532 96380 62534
rect 96436 62532 96460 62534
rect 96516 62532 96540 62534
rect 96596 62532 96620 62534
rect 96676 62532 96682 62534
rect 96374 62523 96682 62532
rect 96896 62280 96948 62286
rect 96896 62222 96948 62228
rect 96374 61500 96682 61509
rect 96374 61498 96380 61500
rect 96436 61498 96460 61500
rect 96516 61498 96540 61500
rect 96596 61498 96620 61500
rect 96676 61498 96682 61500
rect 96436 61446 96438 61498
rect 96618 61446 96620 61498
rect 96374 61444 96380 61446
rect 96436 61444 96460 61446
rect 96516 61444 96540 61446
rect 96596 61444 96620 61446
rect 96676 61444 96682 61446
rect 96374 61435 96682 61444
rect 96252 61396 96304 61402
rect 96252 61338 96304 61344
rect 96908 61266 96936 62222
rect 100392 62144 100444 62150
rect 100392 62086 100444 62092
rect 97034 62044 97342 62053
rect 97034 62042 97040 62044
rect 97096 62042 97120 62044
rect 97176 62042 97200 62044
rect 97256 62042 97280 62044
rect 97336 62042 97342 62044
rect 97096 61990 97098 62042
rect 97278 61990 97280 62042
rect 97034 61988 97040 61990
rect 97096 61988 97120 61990
rect 97176 61988 97200 61990
rect 97256 61988 97280 61990
rect 97336 61988 97342 61990
rect 97034 61979 97342 61988
rect 100404 61985 100432 62086
rect 100390 61976 100446 61985
rect 100390 61911 100446 61920
rect 100208 61804 100260 61810
rect 100208 61746 100260 61752
rect 96896 61260 96948 61266
rect 96896 61202 96948 61208
rect 83924 61192 83976 61198
rect 83924 61134 83976 61140
rect 82452 61124 82504 61130
rect 82452 61066 82504 61072
rect 82820 61124 82872 61130
rect 82820 61066 82872 61072
rect 81716 60784 81768 60790
rect 81716 60726 81768 60732
rect 81532 60648 81584 60654
rect 81532 60590 81584 60596
rect 79508 60512 79560 60518
rect 79508 60454 79560 60460
rect 79692 60512 79744 60518
rect 79692 60454 79744 60460
rect 81440 60512 81492 60518
rect 81440 60454 81492 60460
rect 79232 60104 79284 60110
rect 79232 60046 79284 60052
rect 79520 58721 79548 60454
rect 81348 60104 81400 60110
rect 81348 60046 81400 60052
rect 81360 58750 81388 60046
rect 81452 60042 81480 60454
rect 81728 60314 81756 60726
rect 81808 60648 81860 60654
rect 81808 60590 81860 60596
rect 81716 60308 81768 60314
rect 81716 60250 81768 60256
rect 81440 60036 81492 60042
rect 81440 59978 81492 59984
rect 81348 58744 81400 58750
rect 79506 58712 79562 58721
rect 81348 58686 81400 58692
rect 79506 58647 79562 58656
rect 79138 58576 79194 58585
rect 79138 58511 79194 58520
rect 29182 58168 29238 58177
rect 29182 58103 29238 58112
rect 81820 57905 81848 60590
rect 82832 60314 82860 61066
rect 83832 61056 83884 61062
rect 83832 60998 83884 61004
rect 83844 60858 83872 60998
rect 83832 60852 83884 60858
rect 83832 60794 83884 60800
rect 83936 60738 83964 61134
rect 84016 61056 84068 61062
rect 84016 60998 84068 61004
rect 84028 60790 84056 60998
rect 97034 60956 97342 60965
rect 97034 60954 97040 60956
rect 97096 60954 97120 60956
rect 97176 60954 97200 60956
rect 97256 60954 97280 60956
rect 97336 60954 97342 60956
rect 97096 60902 97098 60954
rect 97278 60902 97280 60954
rect 97034 60900 97040 60902
rect 97096 60900 97120 60902
rect 97176 60900 97200 60902
rect 97256 60900 97280 60902
rect 97336 60900 97342 60902
rect 97034 60891 97342 60900
rect 83844 60710 83964 60738
rect 84016 60784 84068 60790
rect 84016 60726 84068 60732
rect 85580 60784 85632 60790
rect 85580 60726 85632 60732
rect 83280 60512 83332 60518
rect 83280 60454 83332 60460
rect 82820 60308 82872 60314
rect 82820 60250 82872 60256
rect 83292 60246 83320 60454
rect 83280 60240 83332 60246
rect 83280 60182 83332 60188
rect 83844 60110 83872 60710
rect 83924 60648 83976 60654
rect 83924 60590 83976 60596
rect 83936 60178 83964 60590
rect 85592 60314 85620 60726
rect 85672 60648 85724 60654
rect 85672 60590 85724 60596
rect 87604 60648 87656 60654
rect 87604 60590 87656 60596
rect 87880 60648 87932 60654
rect 87880 60590 87932 60596
rect 85684 60314 85712 60590
rect 86132 60512 86184 60518
rect 86132 60454 86184 60460
rect 85580 60308 85632 60314
rect 85580 60250 85632 60256
rect 85672 60308 85724 60314
rect 85672 60250 85724 60256
rect 83924 60172 83976 60178
rect 83924 60114 83976 60120
rect 83832 60104 83884 60110
rect 83832 60046 83884 60052
rect 83936 58041 83964 60114
rect 86144 60110 86172 60454
rect 87616 60314 87644 60590
rect 87892 60518 87920 60590
rect 87880 60512 87932 60518
rect 87880 60454 87932 60460
rect 87604 60308 87656 60314
rect 87604 60250 87656 60256
rect 84384 60104 84436 60110
rect 84384 60046 84436 60052
rect 86132 60104 86184 60110
rect 86132 60046 86184 60052
rect 84396 58818 84424 60046
rect 84384 58812 84436 58818
rect 84384 58754 84436 58760
rect 86144 58585 86172 60046
rect 86130 58576 86186 58585
rect 86130 58511 86186 58520
rect 86144 58177 86172 58511
rect 86130 58168 86186 58177
rect 86130 58103 86186 58112
rect 83922 58032 83978 58041
rect 83922 57967 83978 57976
rect 87892 57905 87920 60454
rect 96374 60412 96682 60421
rect 96374 60410 96380 60412
rect 96436 60410 96460 60412
rect 96516 60410 96540 60412
rect 96596 60410 96620 60412
rect 96676 60410 96682 60412
rect 96436 60358 96438 60410
rect 96618 60358 96620 60410
rect 96374 60356 96380 60358
rect 96436 60356 96460 60358
rect 96516 60356 96540 60358
rect 96596 60356 96620 60358
rect 96676 60356 96682 60358
rect 96374 60347 96682 60356
rect 98930 60412 99238 60421
rect 98930 60410 98936 60412
rect 98992 60410 99016 60412
rect 99072 60410 99096 60412
rect 99152 60410 99176 60412
rect 99232 60410 99238 60412
rect 98992 60358 98994 60410
rect 99174 60358 99176 60410
rect 98930 60356 98936 60358
rect 98992 60356 99016 60358
rect 99072 60356 99096 60358
rect 99152 60356 99176 60358
rect 99232 60356 99238 60358
rect 98930 60347 99238 60356
rect 100220 60314 100248 61746
rect 100392 61600 100444 61606
rect 100392 61542 100444 61548
rect 100404 61305 100432 61542
rect 100390 61296 100446 61305
rect 100390 61231 100446 61240
rect 100390 60616 100446 60625
rect 100390 60551 100392 60560
rect 100444 60551 100446 60560
rect 100392 60522 100444 60528
rect 100208 60308 100260 60314
rect 100208 60250 100260 60256
rect 91744 60240 91796 60246
rect 91744 60182 91796 60188
rect 89536 60104 89588 60110
rect 89720 60104 89772 60110
rect 89588 60052 89720 60058
rect 89536 60046 89772 60052
rect 89548 60030 89760 60046
rect 91756 60042 91784 60182
rect 98368 60104 98420 60110
rect 98368 60046 98420 60052
rect 91744 60036 91796 60042
rect 91744 59978 91796 59984
rect 97034 59868 97342 59877
rect 97034 59866 97040 59868
rect 97096 59866 97120 59868
rect 97176 59866 97200 59868
rect 97256 59866 97280 59868
rect 97336 59866 97342 59868
rect 97096 59814 97098 59866
rect 97278 59814 97280 59866
rect 97034 59812 97040 59814
rect 97096 59812 97120 59814
rect 97176 59812 97200 59814
rect 97256 59812 97280 59814
rect 97336 59812 97342 59814
rect 97034 59803 97342 59812
rect 97356 58812 97408 58818
rect 97356 58754 97408 58760
rect 97264 58676 97316 58682
rect 97264 58618 97316 58624
rect 28170 57896 28226 57905
rect 28170 57831 28226 57840
rect 81806 57896 81862 57905
rect 81806 57831 81862 57840
rect 87878 57896 87934 57905
rect 87878 57831 87934 57840
rect 97080 53984 97132 53990
rect 97080 53926 97132 53932
rect 97092 53825 97120 53926
rect 97078 53816 97134 53825
rect 97078 53751 97134 53760
rect 97276 4185 97304 58618
rect 97368 27606 97396 58754
rect 97448 58744 97500 58750
rect 97448 58686 97500 58692
rect 97460 43314 97488 58686
rect 98274 58576 98330 58585
rect 98274 58511 98330 58520
rect 98288 45966 98316 58511
rect 98380 45966 98408 60046
rect 100392 59968 100444 59974
rect 100390 59936 100392 59945
rect 100444 59936 100446 59945
rect 99666 59868 99974 59877
rect 100390 59871 100446 59880
rect 99666 59866 99672 59868
rect 99728 59866 99752 59868
rect 99808 59866 99832 59868
rect 99888 59866 99912 59868
rect 99968 59866 99974 59868
rect 99728 59814 99730 59866
rect 99910 59814 99912 59866
rect 99666 59812 99672 59814
rect 99728 59812 99752 59814
rect 99808 59812 99832 59814
rect 99888 59812 99912 59814
rect 99968 59812 99974 59814
rect 99666 59803 99974 59812
rect 98930 59324 99238 59333
rect 98930 59322 98936 59324
rect 98992 59322 99016 59324
rect 99072 59322 99096 59324
rect 99152 59322 99176 59324
rect 99232 59322 99238 59324
rect 98992 59270 98994 59322
rect 99174 59270 99176 59322
rect 98930 59268 98936 59270
rect 98992 59268 99016 59270
rect 99072 59268 99096 59270
rect 99152 59268 99176 59270
rect 99232 59268 99238 59270
rect 98930 59259 99238 59268
rect 99666 58780 99974 58789
rect 99666 58778 99672 58780
rect 99728 58778 99752 58780
rect 99808 58778 99832 58780
rect 99888 58778 99912 58780
rect 99968 58778 99974 58780
rect 99728 58726 99730 58778
rect 99910 58726 99912 58778
rect 99666 58724 99672 58726
rect 99728 58724 99752 58726
rect 99808 58724 99832 58726
rect 99888 58724 99912 58726
rect 99968 58724 99974 58726
rect 99666 58715 99974 58724
rect 98930 58236 99238 58245
rect 98930 58234 98936 58236
rect 98992 58234 99016 58236
rect 99072 58234 99096 58236
rect 99152 58234 99176 58236
rect 99232 58234 99238 58236
rect 98992 58182 98994 58234
rect 99174 58182 99176 58234
rect 98930 58180 98936 58182
rect 98992 58180 99016 58182
rect 99072 58180 99096 58182
rect 99152 58180 99176 58182
rect 99232 58180 99238 58182
rect 98930 58171 99238 58180
rect 100114 57896 100170 57905
rect 100114 57831 100170 57840
rect 99666 57692 99974 57701
rect 99666 57690 99672 57692
rect 99728 57690 99752 57692
rect 99808 57690 99832 57692
rect 99888 57690 99912 57692
rect 99968 57690 99974 57692
rect 99728 57638 99730 57690
rect 99910 57638 99912 57690
rect 99666 57636 99672 57638
rect 99728 57636 99752 57638
rect 99808 57636 99832 57638
rect 99888 57636 99912 57638
rect 99968 57636 99974 57638
rect 99666 57627 99974 57636
rect 98930 57148 99238 57157
rect 98930 57146 98936 57148
rect 98992 57146 99016 57148
rect 99072 57146 99096 57148
rect 99152 57146 99176 57148
rect 99232 57146 99238 57148
rect 98992 57094 98994 57146
rect 99174 57094 99176 57146
rect 98930 57092 98936 57094
rect 98992 57092 99016 57094
rect 99072 57092 99096 57094
rect 99152 57092 99176 57094
rect 99232 57092 99238 57094
rect 98930 57083 99238 57092
rect 99666 56604 99974 56613
rect 99666 56602 99672 56604
rect 99728 56602 99752 56604
rect 99808 56602 99832 56604
rect 99888 56602 99912 56604
rect 99968 56602 99974 56604
rect 99728 56550 99730 56602
rect 99910 56550 99912 56602
rect 99666 56548 99672 56550
rect 99728 56548 99752 56550
rect 99808 56548 99832 56550
rect 99888 56548 99912 56550
rect 99968 56548 99974 56550
rect 99666 56539 99974 56548
rect 98930 56060 99238 56069
rect 98930 56058 98936 56060
rect 98992 56058 99016 56060
rect 99072 56058 99096 56060
rect 99152 56058 99176 56060
rect 99232 56058 99238 56060
rect 98992 56006 98994 56058
rect 99174 56006 99176 56058
rect 98930 56004 98936 56006
rect 98992 56004 99016 56006
rect 99072 56004 99096 56006
rect 99152 56004 99176 56006
rect 99232 56004 99238 56006
rect 98930 55995 99238 56004
rect 99666 55516 99974 55525
rect 99666 55514 99672 55516
rect 99728 55514 99752 55516
rect 99808 55514 99832 55516
rect 99888 55514 99912 55516
rect 99968 55514 99974 55516
rect 99728 55462 99730 55514
rect 99910 55462 99912 55514
rect 99666 55460 99672 55462
rect 99728 55460 99752 55462
rect 99808 55460 99832 55462
rect 99888 55460 99912 55462
rect 99968 55460 99974 55462
rect 99666 55451 99974 55460
rect 98930 54972 99238 54981
rect 98930 54970 98936 54972
rect 98992 54970 99016 54972
rect 99072 54970 99096 54972
rect 99152 54970 99176 54972
rect 99232 54970 99238 54972
rect 98992 54918 98994 54970
rect 99174 54918 99176 54970
rect 98930 54916 98936 54918
rect 98992 54916 99016 54918
rect 99072 54916 99096 54918
rect 99152 54916 99176 54918
rect 99232 54916 99238 54918
rect 98930 54907 99238 54916
rect 99666 54428 99974 54437
rect 99666 54426 99672 54428
rect 99728 54426 99752 54428
rect 99808 54426 99832 54428
rect 99888 54426 99912 54428
rect 99968 54426 99974 54428
rect 99728 54374 99730 54426
rect 99910 54374 99912 54426
rect 99666 54372 99672 54374
rect 99728 54372 99752 54374
rect 99808 54372 99832 54374
rect 99888 54372 99912 54374
rect 99968 54372 99974 54374
rect 99666 54363 99974 54372
rect 98930 53884 99238 53893
rect 98930 53882 98936 53884
rect 98992 53882 99016 53884
rect 99072 53882 99096 53884
rect 99152 53882 99176 53884
rect 99232 53882 99238 53884
rect 98992 53830 98994 53882
rect 99174 53830 99176 53882
rect 98930 53828 98936 53830
rect 98992 53828 99016 53830
rect 99072 53828 99096 53830
rect 99152 53828 99176 53830
rect 99232 53828 99238 53830
rect 98930 53819 99238 53828
rect 99666 53340 99974 53349
rect 99666 53338 99672 53340
rect 99728 53338 99752 53340
rect 99808 53338 99832 53340
rect 99888 53338 99912 53340
rect 99968 53338 99974 53340
rect 99728 53286 99730 53338
rect 99910 53286 99912 53338
rect 99666 53284 99672 53286
rect 99728 53284 99752 53286
rect 99808 53284 99832 53286
rect 99888 53284 99912 53286
rect 99968 53284 99974 53286
rect 99666 53275 99974 53284
rect 98930 52796 99238 52805
rect 98930 52794 98936 52796
rect 98992 52794 99016 52796
rect 99072 52794 99096 52796
rect 99152 52794 99176 52796
rect 99232 52794 99238 52796
rect 98992 52742 98994 52794
rect 99174 52742 99176 52794
rect 98930 52740 98936 52742
rect 98992 52740 99016 52742
rect 99072 52740 99096 52742
rect 99152 52740 99176 52742
rect 99232 52740 99238 52742
rect 98930 52731 99238 52740
rect 99666 52252 99974 52261
rect 99666 52250 99672 52252
rect 99728 52250 99752 52252
rect 99808 52250 99832 52252
rect 99888 52250 99912 52252
rect 99968 52250 99974 52252
rect 99728 52198 99730 52250
rect 99910 52198 99912 52250
rect 99666 52196 99672 52198
rect 99728 52196 99752 52198
rect 99808 52196 99832 52198
rect 99888 52196 99912 52198
rect 99968 52196 99974 52198
rect 99666 52187 99974 52196
rect 98930 51708 99238 51717
rect 98930 51706 98936 51708
rect 98992 51706 99016 51708
rect 99072 51706 99096 51708
rect 99152 51706 99176 51708
rect 99232 51706 99238 51708
rect 98992 51654 98994 51706
rect 99174 51654 99176 51706
rect 98930 51652 98936 51654
rect 98992 51652 99016 51654
rect 99072 51652 99096 51654
rect 99152 51652 99176 51654
rect 99232 51652 99238 51654
rect 98930 51643 99238 51652
rect 99666 51164 99974 51173
rect 99666 51162 99672 51164
rect 99728 51162 99752 51164
rect 99808 51162 99832 51164
rect 99888 51162 99912 51164
rect 99968 51162 99974 51164
rect 99728 51110 99730 51162
rect 99910 51110 99912 51162
rect 99666 51108 99672 51110
rect 99728 51108 99752 51110
rect 99808 51108 99832 51110
rect 99888 51108 99912 51110
rect 99968 51108 99974 51110
rect 99666 51099 99974 51108
rect 98930 50620 99238 50629
rect 98930 50618 98936 50620
rect 98992 50618 99016 50620
rect 99072 50618 99096 50620
rect 99152 50618 99176 50620
rect 99232 50618 99238 50620
rect 98992 50566 98994 50618
rect 99174 50566 99176 50618
rect 98930 50564 98936 50566
rect 98992 50564 99016 50566
rect 99072 50564 99096 50566
rect 99152 50564 99176 50566
rect 99232 50564 99238 50566
rect 98930 50555 99238 50564
rect 99666 50076 99974 50085
rect 99666 50074 99672 50076
rect 99728 50074 99752 50076
rect 99808 50074 99832 50076
rect 99888 50074 99912 50076
rect 99968 50074 99974 50076
rect 99728 50022 99730 50074
rect 99910 50022 99912 50074
rect 99666 50020 99672 50022
rect 99728 50020 99752 50022
rect 99808 50020 99832 50022
rect 99888 50020 99912 50022
rect 99968 50020 99974 50022
rect 99666 50011 99974 50020
rect 98930 49532 99238 49541
rect 98930 49530 98936 49532
rect 98992 49530 99016 49532
rect 99072 49530 99096 49532
rect 99152 49530 99176 49532
rect 99232 49530 99238 49532
rect 98992 49478 98994 49530
rect 99174 49478 99176 49530
rect 98930 49476 98936 49478
rect 98992 49476 99016 49478
rect 99072 49476 99096 49478
rect 99152 49476 99176 49478
rect 99232 49476 99238 49478
rect 98930 49467 99238 49476
rect 99666 48988 99974 48997
rect 99666 48986 99672 48988
rect 99728 48986 99752 48988
rect 99808 48986 99832 48988
rect 99888 48986 99912 48988
rect 99968 48986 99974 48988
rect 99728 48934 99730 48986
rect 99910 48934 99912 48986
rect 99666 48932 99672 48934
rect 99728 48932 99752 48934
rect 99808 48932 99832 48934
rect 99888 48932 99912 48934
rect 99968 48932 99974 48934
rect 99666 48923 99974 48932
rect 98930 48444 99238 48453
rect 98930 48442 98936 48444
rect 98992 48442 99016 48444
rect 99072 48442 99096 48444
rect 99152 48442 99176 48444
rect 99232 48442 99238 48444
rect 98992 48390 98994 48442
rect 99174 48390 99176 48442
rect 98930 48388 98936 48390
rect 98992 48388 99016 48390
rect 99072 48388 99096 48390
rect 99152 48388 99176 48390
rect 99232 48388 99238 48390
rect 98930 48379 99238 48388
rect 99666 47900 99974 47909
rect 99666 47898 99672 47900
rect 99728 47898 99752 47900
rect 99808 47898 99832 47900
rect 99888 47898 99912 47900
rect 99968 47898 99974 47900
rect 99728 47846 99730 47898
rect 99910 47846 99912 47898
rect 99666 47844 99672 47846
rect 99728 47844 99752 47846
rect 99808 47844 99832 47846
rect 99888 47844 99912 47846
rect 99968 47844 99974 47846
rect 99666 47835 99974 47844
rect 98930 47356 99238 47365
rect 98930 47354 98936 47356
rect 98992 47354 99016 47356
rect 99072 47354 99096 47356
rect 99152 47354 99176 47356
rect 99232 47354 99238 47356
rect 98992 47302 98994 47354
rect 99174 47302 99176 47354
rect 98930 47300 98936 47302
rect 98992 47300 99016 47302
rect 99072 47300 99096 47302
rect 99152 47300 99176 47302
rect 99232 47300 99238 47302
rect 98930 47291 99238 47300
rect 99666 46812 99974 46821
rect 99666 46810 99672 46812
rect 99728 46810 99752 46812
rect 99808 46810 99832 46812
rect 99888 46810 99912 46812
rect 99968 46810 99974 46812
rect 99728 46758 99730 46810
rect 99910 46758 99912 46810
rect 99666 46756 99672 46758
rect 99728 46756 99752 46758
rect 99808 46756 99832 46758
rect 99888 46756 99912 46758
rect 99968 46756 99974 46758
rect 99666 46747 99974 46756
rect 98930 46268 99238 46277
rect 98930 46266 98936 46268
rect 98992 46266 99016 46268
rect 99072 46266 99096 46268
rect 99152 46266 99176 46268
rect 99232 46266 99238 46268
rect 98992 46214 98994 46266
rect 99174 46214 99176 46266
rect 98930 46212 98936 46214
rect 98992 46212 99016 46214
rect 99072 46212 99096 46214
rect 99152 46212 99176 46214
rect 99232 46212 99238 46214
rect 98930 46203 99238 46212
rect 98552 46096 98604 46102
rect 98552 46038 98604 46044
rect 98276 45960 98328 45966
rect 98276 45902 98328 45908
rect 98368 45960 98420 45966
rect 98368 45902 98420 45908
rect 98184 45892 98236 45898
rect 98184 45834 98236 45840
rect 98196 44742 98224 45834
rect 98288 45082 98316 45902
rect 98276 45076 98328 45082
rect 98276 45018 98328 45024
rect 98380 44810 98408 45902
rect 98368 44804 98420 44810
rect 98368 44746 98420 44752
rect 98184 44736 98236 44742
rect 98184 44678 98236 44684
rect 97448 43308 97500 43314
rect 97448 43250 97500 43256
rect 98196 40934 98224 44678
rect 98276 43308 98328 43314
rect 98276 43250 98328 43256
rect 98184 40928 98236 40934
rect 98184 40870 98236 40876
rect 97356 27600 97408 27606
rect 97356 27542 97408 27548
rect 98092 25152 98144 25158
rect 98092 25094 98144 25100
rect 98104 23526 98132 25094
rect 98092 23520 98144 23526
rect 98092 23462 98144 23468
rect 97356 22772 97408 22778
rect 97356 22714 97408 22720
rect 97262 4176 97318 4185
rect 97262 4111 97318 4120
rect 2686 3904 2742 3913
rect 1312 3836 1448 3845
rect 2686 3839 2742 3848
rect 1368 3834 1392 3836
rect 1374 3782 1386 3834
rect 1368 3780 1392 3782
rect 1312 3771 1448 3780
rect 97368 3641 97396 22714
rect 97540 21956 97592 21962
rect 97540 21898 97592 21904
rect 97552 3777 97580 21898
rect 98196 19145 98224 40870
rect 98288 35698 98316 43250
rect 98368 43104 98420 43110
rect 98368 43046 98420 43052
rect 98380 41206 98408 43046
rect 98368 41200 98420 41206
rect 98368 41142 98420 41148
rect 98460 41064 98512 41070
rect 98460 41006 98512 41012
rect 98472 40730 98500 41006
rect 98460 40724 98512 40730
rect 98460 40666 98512 40672
rect 98564 40526 98592 46038
rect 99666 45724 99974 45733
rect 99666 45722 99672 45724
rect 99728 45722 99752 45724
rect 99808 45722 99832 45724
rect 99888 45722 99912 45724
rect 99968 45722 99974 45724
rect 99728 45670 99730 45722
rect 99910 45670 99912 45722
rect 99666 45668 99672 45670
rect 99728 45668 99752 45670
rect 99808 45668 99832 45670
rect 99888 45668 99912 45670
rect 99968 45668 99974 45670
rect 99666 45659 99974 45668
rect 98930 45180 99238 45189
rect 98930 45178 98936 45180
rect 98992 45178 99016 45180
rect 99072 45178 99096 45180
rect 99152 45178 99176 45180
rect 99232 45178 99238 45180
rect 98992 45126 98994 45178
rect 99174 45126 99176 45178
rect 98930 45124 98936 45126
rect 98992 45124 99016 45126
rect 99072 45124 99096 45126
rect 99152 45124 99176 45126
rect 99232 45124 99238 45126
rect 98930 45115 99238 45124
rect 98644 44736 98696 44742
rect 98644 44678 98696 44684
rect 98552 40520 98604 40526
rect 98552 40462 98604 40468
rect 98656 40458 98684 44678
rect 99666 44636 99974 44645
rect 99666 44634 99672 44636
rect 99728 44634 99752 44636
rect 99808 44634 99832 44636
rect 99888 44634 99912 44636
rect 99968 44634 99974 44636
rect 99728 44582 99730 44634
rect 99910 44582 99912 44634
rect 99666 44580 99672 44582
rect 99728 44580 99752 44582
rect 99808 44580 99832 44582
rect 99888 44580 99912 44582
rect 99968 44580 99974 44582
rect 99666 44571 99974 44580
rect 98930 44092 99238 44101
rect 98930 44090 98936 44092
rect 98992 44090 99016 44092
rect 99072 44090 99096 44092
rect 99152 44090 99176 44092
rect 99232 44090 99238 44092
rect 98992 44038 98994 44090
rect 99174 44038 99176 44090
rect 98930 44036 98936 44038
rect 98992 44036 99016 44038
rect 99072 44036 99096 44038
rect 99152 44036 99176 44038
rect 99232 44036 99238 44038
rect 98930 44027 99238 44036
rect 99666 43548 99974 43557
rect 99666 43546 99672 43548
rect 99728 43546 99752 43548
rect 99808 43546 99832 43548
rect 99888 43546 99912 43548
rect 99968 43546 99974 43548
rect 99728 43494 99730 43546
rect 99910 43494 99912 43546
rect 99666 43492 99672 43494
rect 99728 43492 99752 43494
rect 99808 43492 99832 43494
rect 99888 43492 99912 43494
rect 99968 43492 99974 43494
rect 99666 43483 99974 43492
rect 98930 43004 99238 43013
rect 98930 43002 98936 43004
rect 98992 43002 99016 43004
rect 99072 43002 99096 43004
rect 99152 43002 99176 43004
rect 99232 43002 99238 43004
rect 98992 42950 98994 43002
rect 99174 42950 99176 43002
rect 98930 42948 98936 42950
rect 98992 42948 99016 42950
rect 99072 42948 99096 42950
rect 99152 42948 99176 42950
rect 99232 42948 99238 42950
rect 98930 42939 99238 42948
rect 99666 42460 99974 42469
rect 99666 42458 99672 42460
rect 99728 42458 99752 42460
rect 99808 42458 99832 42460
rect 99888 42458 99912 42460
rect 99968 42458 99974 42460
rect 99728 42406 99730 42458
rect 99910 42406 99912 42458
rect 99666 42404 99672 42406
rect 99728 42404 99752 42406
rect 99808 42404 99832 42406
rect 99888 42404 99912 42406
rect 99968 42404 99974 42406
rect 99666 42395 99974 42404
rect 98930 41916 99238 41925
rect 98930 41914 98936 41916
rect 98992 41914 99016 41916
rect 99072 41914 99096 41916
rect 99152 41914 99176 41916
rect 99232 41914 99238 41916
rect 98992 41862 98994 41914
rect 99174 41862 99176 41914
rect 98930 41860 98936 41862
rect 98992 41860 99016 41862
rect 99072 41860 99096 41862
rect 99152 41860 99176 41862
rect 99232 41860 99238 41862
rect 98930 41851 99238 41860
rect 99666 41372 99974 41381
rect 99666 41370 99672 41372
rect 99728 41370 99752 41372
rect 99808 41370 99832 41372
rect 99888 41370 99912 41372
rect 99968 41370 99974 41372
rect 99728 41318 99730 41370
rect 99910 41318 99912 41370
rect 99666 41316 99672 41318
rect 99728 41316 99752 41318
rect 99808 41316 99832 41318
rect 99888 41316 99912 41318
rect 99968 41316 99974 41318
rect 99666 41307 99974 41316
rect 100128 41070 100156 57831
rect 100116 41064 100168 41070
rect 100116 41006 100168 41012
rect 98930 40828 99238 40837
rect 98930 40826 98936 40828
rect 98992 40826 99016 40828
rect 99072 40826 99096 40828
rect 99152 40826 99176 40828
rect 99232 40826 99238 40828
rect 98992 40774 98994 40826
rect 99174 40774 99176 40826
rect 98930 40772 98936 40774
rect 98992 40772 99016 40774
rect 99072 40772 99096 40774
rect 99152 40772 99176 40774
rect 99232 40772 99238 40774
rect 98930 40763 99238 40772
rect 98644 40452 98696 40458
rect 98644 40394 98696 40400
rect 99666 40284 99974 40293
rect 99666 40282 99672 40284
rect 99728 40282 99752 40284
rect 99808 40282 99832 40284
rect 99888 40282 99912 40284
rect 99968 40282 99974 40284
rect 99728 40230 99730 40282
rect 99910 40230 99912 40282
rect 99666 40228 99672 40230
rect 99728 40228 99752 40230
rect 99808 40228 99832 40230
rect 99888 40228 99912 40230
rect 99968 40228 99974 40230
rect 99666 40219 99974 40228
rect 98930 39740 99238 39749
rect 98930 39738 98936 39740
rect 98992 39738 99016 39740
rect 99072 39738 99096 39740
rect 99152 39738 99176 39740
rect 99232 39738 99238 39740
rect 98992 39686 98994 39738
rect 99174 39686 99176 39738
rect 98930 39684 98936 39686
rect 98992 39684 99016 39686
rect 99072 39684 99096 39686
rect 99152 39684 99176 39686
rect 99232 39684 99238 39686
rect 98930 39675 99238 39684
rect 99666 39196 99974 39205
rect 99666 39194 99672 39196
rect 99728 39194 99752 39196
rect 99808 39194 99832 39196
rect 99888 39194 99912 39196
rect 99968 39194 99974 39196
rect 99728 39142 99730 39194
rect 99910 39142 99912 39194
rect 99666 39140 99672 39142
rect 99728 39140 99752 39142
rect 99808 39140 99832 39142
rect 99888 39140 99912 39142
rect 99968 39140 99974 39142
rect 99666 39131 99974 39140
rect 98930 38652 99238 38661
rect 98930 38650 98936 38652
rect 98992 38650 99016 38652
rect 99072 38650 99096 38652
rect 99152 38650 99176 38652
rect 99232 38650 99238 38652
rect 98992 38598 98994 38650
rect 99174 38598 99176 38650
rect 98930 38596 98936 38598
rect 98992 38596 99016 38598
rect 99072 38596 99096 38598
rect 99152 38596 99176 38598
rect 99232 38596 99238 38598
rect 98930 38587 99238 38596
rect 99666 38108 99974 38117
rect 99666 38106 99672 38108
rect 99728 38106 99752 38108
rect 99808 38106 99832 38108
rect 99888 38106 99912 38108
rect 99968 38106 99974 38108
rect 99728 38054 99730 38106
rect 99910 38054 99912 38106
rect 99666 38052 99672 38054
rect 99728 38052 99752 38054
rect 99808 38052 99832 38054
rect 99888 38052 99912 38054
rect 99968 38052 99974 38054
rect 99666 38043 99974 38052
rect 98930 37564 99238 37573
rect 98930 37562 98936 37564
rect 98992 37562 99016 37564
rect 99072 37562 99096 37564
rect 99152 37562 99176 37564
rect 99232 37562 99238 37564
rect 98992 37510 98994 37562
rect 99174 37510 99176 37562
rect 98930 37508 98936 37510
rect 98992 37508 99016 37510
rect 99072 37508 99096 37510
rect 99152 37508 99176 37510
rect 99232 37508 99238 37510
rect 98930 37499 99238 37508
rect 99666 37020 99974 37029
rect 99666 37018 99672 37020
rect 99728 37018 99752 37020
rect 99808 37018 99832 37020
rect 99888 37018 99912 37020
rect 99968 37018 99974 37020
rect 99728 36966 99730 37018
rect 99910 36966 99912 37018
rect 99666 36964 99672 36966
rect 99728 36964 99752 36966
rect 99808 36964 99832 36966
rect 99888 36964 99912 36966
rect 99968 36964 99974 36966
rect 99666 36955 99974 36964
rect 98930 36476 99238 36485
rect 98930 36474 98936 36476
rect 98992 36474 99016 36476
rect 99072 36474 99096 36476
rect 99152 36474 99176 36476
rect 99232 36474 99238 36476
rect 98992 36422 98994 36474
rect 99174 36422 99176 36474
rect 98930 36420 98936 36422
rect 98992 36420 99016 36422
rect 99072 36420 99096 36422
rect 99152 36420 99176 36422
rect 99232 36420 99238 36422
rect 98930 36411 99238 36420
rect 99666 35932 99974 35941
rect 99666 35930 99672 35932
rect 99728 35930 99752 35932
rect 99808 35930 99832 35932
rect 99888 35930 99912 35932
rect 99968 35930 99974 35932
rect 99728 35878 99730 35930
rect 99910 35878 99912 35930
rect 99666 35876 99672 35878
rect 99728 35876 99752 35878
rect 99808 35876 99832 35878
rect 99888 35876 99912 35878
rect 99968 35876 99974 35878
rect 99666 35867 99974 35876
rect 98276 35692 98328 35698
rect 98276 35634 98328 35640
rect 98460 35692 98512 35698
rect 98460 35634 98512 35640
rect 98472 34610 98500 35634
rect 98736 35488 98788 35494
rect 98736 35430 98788 35436
rect 98460 34604 98512 34610
rect 98460 34546 98512 34552
rect 98368 34536 98420 34542
rect 98368 34478 98420 34484
rect 98380 30666 98408 34478
rect 98368 30660 98420 30666
rect 98368 30602 98420 30608
rect 98276 30592 98328 30598
rect 98276 30534 98328 30540
rect 98288 29102 98316 30534
rect 98472 29646 98500 34546
rect 98748 31822 98776 35430
rect 98930 35388 99238 35397
rect 98930 35386 98936 35388
rect 98992 35386 99016 35388
rect 99072 35386 99096 35388
rect 99152 35386 99176 35388
rect 99232 35386 99238 35388
rect 98992 35334 98994 35386
rect 99174 35334 99176 35386
rect 98930 35332 98936 35334
rect 98992 35332 99016 35334
rect 99072 35332 99096 35334
rect 99152 35332 99176 35334
rect 99232 35332 99238 35334
rect 98930 35323 99238 35332
rect 99666 34844 99974 34853
rect 99666 34842 99672 34844
rect 99728 34842 99752 34844
rect 99808 34842 99832 34844
rect 99888 34842 99912 34844
rect 99968 34842 99974 34844
rect 99728 34790 99730 34842
rect 99910 34790 99912 34842
rect 99666 34788 99672 34790
rect 99728 34788 99752 34790
rect 99808 34788 99832 34790
rect 99888 34788 99912 34790
rect 99968 34788 99974 34790
rect 99666 34779 99974 34788
rect 98930 34300 99238 34309
rect 98930 34298 98936 34300
rect 98992 34298 99016 34300
rect 99072 34298 99096 34300
rect 99152 34298 99176 34300
rect 99232 34298 99238 34300
rect 98992 34246 98994 34298
rect 99174 34246 99176 34298
rect 98930 34244 98936 34246
rect 98992 34244 99016 34246
rect 99072 34244 99096 34246
rect 99152 34244 99176 34246
rect 99232 34244 99238 34246
rect 98930 34235 99238 34244
rect 99666 33756 99974 33765
rect 99666 33754 99672 33756
rect 99728 33754 99752 33756
rect 99808 33754 99832 33756
rect 99888 33754 99912 33756
rect 99968 33754 99974 33756
rect 99728 33702 99730 33754
rect 99910 33702 99912 33754
rect 99666 33700 99672 33702
rect 99728 33700 99752 33702
rect 99808 33700 99832 33702
rect 99888 33700 99912 33702
rect 99968 33700 99974 33702
rect 99666 33691 99974 33700
rect 98930 33212 99238 33221
rect 98930 33210 98936 33212
rect 98992 33210 99016 33212
rect 99072 33210 99096 33212
rect 99152 33210 99176 33212
rect 99232 33210 99238 33212
rect 98992 33158 98994 33210
rect 99174 33158 99176 33210
rect 98930 33156 98936 33158
rect 98992 33156 99016 33158
rect 99072 33156 99096 33158
rect 99152 33156 99176 33158
rect 99232 33156 99238 33158
rect 98930 33147 99238 33156
rect 99666 32668 99974 32677
rect 99666 32666 99672 32668
rect 99728 32666 99752 32668
rect 99808 32666 99832 32668
rect 99888 32666 99912 32668
rect 99968 32666 99974 32668
rect 99728 32614 99730 32666
rect 99910 32614 99912 32666
rect 99666 32612 99672 32614
rect 99728 32612 99752 32614
rect 99808 32612 99832 32614
rect 99888 32612 99912 32614
rect 99968 32612 99974 32614
rect 99666 32603 99974 32612
rect 98930 32124 99238 32133
rect 98930 32122 98936 32124
rect 98992 32122 99016 32124
rect 99072 32122 99096 32124
rect 99152 32122 99176 32124
rect 99232 32122 99238 32124
rect 98992 32070 98994 32122
rect 99174 32070 99176 32122
rect 98930 32068 98936 32070
rect 98992 32068 99016 32070
rect 99072 32068 99096 32070
rect 99152 32068 99176 32070
rect 99232 32068 99238 32070
rect 98930 32059 99238 32068
rect 100128 31906 100156 41006
rect 100208 40452 100260 40458
rect 100208 40394 100260 40400
rect 100220 35894 100248 40394
rect 100220 35866 100340 35894
rect 99380 31884 99432 31890
rect 99380 31826 99432 31832
rect 99840 31884 99892 31890
rect 100128 31878 100248 31906
rect 99840 31826 99892 31832
rect 98736 31816 98788 31822
rect 98736 31758 98788 31764
rect 98930 31036 99238 31045
rect 98930 31034 98936 31036
rect 98992 31034 99016 31036
rect 99072 31034 99096 31036
rect 99152 31034 99176 31036
rect 99232 31034 99238 31036
rect 98992 30982 98994 31034
rect 99174 30982 99176 31034
rect 98930 30980 98936 30982
rect 98992 30980 99016 30982
rect 99072 30980 99096 30982
rect 99152 30980 99176 30982
rect 99232 30980 99238 30982
rect 98930 30971 99238 30980
rect 99392 30258 99420 31826
rect 99852 31770 99880 31826
rect 100220 31822 100248 31878
rect 100208 31816 100260 31822
rect 99852 31742 100064 31770
rect 100208 31758 100260 31764
rect 99666 31580 99974 31589
rect 99666 31578 99672 31580
rect 99728 31578 99752 31580
rect 99808 31578 99832 31580
rect 99888 31578 99912 31580
rect 99968 31578 99974 31580
rect 99728 31526 99730 31578
rect 99910 31526 99912 31578
rect 99666 31524 99672 31526
rect 99728 31524 99752 31526
rect 99808 31524 99832 31526
rect 99888 31524 99912 31526
rect 99968 31524 99974 31526
rect 99666 31515 99974 31524
rect 99564 30592 99616 30598
rect 99564 30534 99616 30540
rect 99380 30252 99432 30258
rect 99380 30194 99432 30200
rect 99380 30048 99432 30054
rect 99380 29990 99432 29996
rect 98930 29948 99238 29957
rect 98930 29946 98936 29948
rect 98992 29946 99016 29948
rect 99072 29946 99096 29948
rect 99152 29946 99176 29948
rect 99232 29946 99238 29948
rect 98992 29894 98994 29946
rect 99174 29894 99176 29946
rect 98930 29892 98936 29894
rect 98992 29892 99016 29894
rect 99072 29892 99096 29894
rect 99152 29892 99176 29894
rect 99232 29892 99238 29894
rect 98930 29883 99238 29892
rect 98460 29640 98512 29646
rect 98460 29582 98512 29588
rect 98736 29640 98788 29646
rect 98736 29582 98788 29588
rect 98644 29504 98696 29510
rect 98644 29446 98696 29452
rect 98276 29096 98328 29102
rect 98276 29038 98328 29044
rect 98552 29028 98604 29034
rect 98552 28970 98604 28976
rect 98368 27600 98420 27606
rect 98368 27542 98420 27548
rect 98380 26450 98408 27542
rect 98368 26444 98420 26450
rect 98368 26386 98420 26392
rect 98380 25974 98408 26386
rect 98368 25968 98420 25974
rect 98368 25910 98420 25916
rect 98368 25832 98420 25838
rect 98368 25774 98420 25780
rect 98276 25696 98328 25702
rect 98276 25638 98328 25644
rect 98288 23730 98316 25638
rect 98380 24206 98408 25774
rect 98564 24818 98592 28970
rect 98656 25362 98684 29446
rect 98748 29170 98776 29582
rect 99392 29170 99420 29990
rect 98736 29164 98788 29170
rect 98736 29106 98788 29112
rect 99380 29164 99432 29170
rect 99380 29106 99432 29112
rect 98748 25838 98776 29106
rect 99288 29096 99340 29102
rect 99288 29038 99340 29044
rect 98930 28860 99238 28869
rect 98930 28858 98936 28860
rect 98992 28858 99016 28860
rect 99072 28858 99096 28860
rect 99152 28858 99176 28860
rect 99232 28858 99238 28860
rect 98992 28806 98994 28858
rect 99174 28806 99176 28858
rect 98930 28804 98936 28806
rect 98992 28804 99016 28806
rect 99072 28804 99096 28806
rect 99152 28804 99176 28806
rect 99232 28804 99238 28806
rect 98930 28795 99238 28804
rect 98930 27772 99238 27781
rect 98930 27770 98936 27772
rect 98992 27770 99016 27772
rect 99072 27770 99096 27772
rect 99152 27770 99176 27772
rect 99232 27770 99238 27772
rect 98992 27718 98994 27770
rect 99174 27718 99176 27770
rect 98930 27716 98936 27718
rect 98992 27716 99016 27718
rect 99072 27716 99096 27718
rect 99152 27716 99176 27718
rect 99232 27716 99238 27718
rect 98930 27707 99238 27716
rect 98930 26684 99238 26693
rect 98930 26682 98936 26684
rect 98992 26682 99016 26684
rect 99072 26682 99096 26684
rect 99152 26682 99176 26684
rect 99232 26682 99238 26684
rect 98992 26630 98994 26682
rect 99174 26630 99176 26682
rect 98930 26628 98936 26630
rect 98992 26628 99016 26630
rect 99072 26628 99096 26630
rect 99152 26628 99176 26630
rect 99232 26628 99238 26630
rect 98930 26619 99238 26628
rect 98736 25832 98788 25838
rect 98736 25774 98788 25780
rect 99300 25770 99328 29038
rect 99472 29028 99524 29034
rect 99472 28970 99524 28976
rect 99484 27470 99512 28970
rect 99576 27606 99604 30534
rect 99666 30492 99974 30501
rect 99666 30490 99672 30492
rect 99728 30490 99752 30492
rect 99808 30490 99832 30492
rect 99888 30490 99912 30492
rect 99968 30490 99974 30492
rect 99728 30438 99730 30490
rect 99910 30438 99912 30490
rect 99666 30436 99672 30438
rect 99728 30436 99752 30438
rect 99808 30436 99832 30438
rect 99888 30436 99912 30438
rect 99968 30436 99974 30438
rect 99666 30427 99974 30436
rect 99666 29404 99974 29413
rect 99666 29402 99672 29404
rect 99728 29402 99752 29404
rect 99808 29402 99832 29404
rect 99888 29402 99912 29404
rect 99968 29402 99974 29404
rect 99728 29350 99730 29402
rect 99910 29350 99912 29402
rect 99666 29348 99672 29350
rect 99728 29348 99752 29350
rect 99808 29348 99832 29350
rect 99888 29348 99912 29350
rect 99968 29348 99974 29350
rect 99666 29339 99974 29348
rect 100036 29034 100064 31742
rect 100220 30734 100248 31758
rect 100208 30728 100260 30734
rect 100208 30670 100260 30676
rect 100116 30252 100168 30258
rect 100116 30194 100168 30200
rect 100024 29028 100076 29034
rect 100024 28970 100076 28976
rect 99666 28316 99974 28325
rect 99666 28314 99672 28316
rect 99728 28314 99752 28316
rect 99808 28314 99832 28316
rect 99888 28314 99912 28316
rect 99968 28314 99974 28316
rect 99728 28262 99730 28314
rect 99910 28262 99912 28314
rect 99666 28260 99672 28262
rect 99728 28260 99752 28262
rect 99808 28260 99832 28262
rect 99888 28260 99912 28262
rect 99968 28260 99974 28262
rect 99666 28251 99974 28260
rect 99564 27600 99616 27606
rect 99564 27542 99616 27548
rect 99472 27464 99524 27470
rect 99472 27406 99524 27412
rect 100024 27464 100076 27470
rect 100024 27406 100076 27412
rect 99564 27396 99616 27402
rect 99564 27338 99616 27344
rect 99576 25906 99604 27338
rect 99666 27228 99974 27237
rect 99666 27226 99672 27228
rect 99728 27226 99752 27228
rect 99808 27226 99832 27228
rect 99888 27226 99912 27228
rect 99968 27226 99974 27228
rect 99728 27174 99730 27226
rect 99910 27174 99912 27226
rect 99666 27172 99672 27174
rect 99728 27172 99752 27174
rect 99808 27172 99832 27174
rect 99888 27172 99912 27174
rect 99968 27172 99974 27174
rect 99666 27163 99974 27172
rect 99666 26140 99974 26149
rect 99666 26138 99672 26140
rect 99728 26138 99752 26140
rect 99808 26138 99832 26140
rect 99888 26138 99912 26140
rect 99968 26138 99974 26140
rect 99728 26086 99730 26138
rect 99910 26086 99912 26138
rect 99666 26084 99672 26086
rect 99728 26084 99752 26086
rect 99808 26084 99832 26086
rect 99888 26084 99912 26086
rect 99968 26084 99974 26086
rect 99666 26075 99974 26084
rect 100036 26042 100064 27406
rect 100128 27402 100156 30194
rect 100116 27396 100168 27402
rect 100116 27338 100168 27344
rect 100024 26036 100076 26042
rect 100024 25978 100076 25984
rect 99564 25900 99616 25906
rect 99564 25842 99616 25848
rect 98828 25764 98880 25770
rect 98828 25706 98880 25712
rect 99288 25764 99340 25770
rect 99288 25706 99340 25712
rect 98644 25356 98696 25362
rect 98644 25298 98696 25304
rect 98552 24812 98604 24818
rect 98552 24754 98604 24760
rect 98552 24608 98604 24614
rect 98552 24550 98604 24556
rect 98368 24200 98420 24206
rect 98368 24142 98420 24148
rect 98460 24064 98512 24070
rect 98460 24006 98512 24012
rect 98276 23724 98328 23730
rect 98276 23666 98328 23672
rect 98368 23520 98420 23526
rect 98368 23462 98420 23468
rect 98380 22778 98408 23462
rect 98368 22772 98420 22778
rect 98368 22714 98420 22720
rect 98276 22568 98328 22574
rect 98276 22510 98328 22516
rect 98288 21962 98316 22510
rect 98276 21956 98328 21962
rect 98276 21898 98328 21904
rect 98472 19786 98500 24006
rect 98564 22574 98592 24550
rect 98736 23860 98788 23866
rect 98736 23802 98788 23808
rect 98748 22778 98776 23802
rect 98736 22772 98788 22778
rect 98736 22714 98788 22720
rect 98552 22568 98604 22574
rect 98552 22510 98604 22516
rect 98552 22432 98604 22438
rect 98552 22374 98604 22380
rect 98460 19780 98512 19786
rect 98460 19722 98512 19728
rect 98368 19712 98420 19718
rect 98368 19654 98420 19660
rect 98380 19310 98408 19654
rect 98368 19304 98420 19310
rect 98368 19246 98420 19252
rect 98182 19136 98238 19145
rect 98182 19071 98238 19080
rect 98380 6914 98408 19246
rect 98460 19168 98512 19174
rect 98460 19110 98512 19116
rect 98472 18290 98500 19110
rect 98460 18284 98512 18290
rect 98460 18226 98512 18232
rect 98564 16289 98592 22374
rect 98748 21962 98776 22714
rect 98840 22438 98868 25706
rect 98930 25596 99238 25605
rect 98930 25594 98936 25596
rect 98992 25594 99016 25596
rect 99072 25594 99096 25596
rect 99152 25594 99176 25596
rect 99232 25594 99238 25596
rect 98992 25542 98994 25594
rect 99174 25542 99176 25594
rect 98930 25540 98936 25542
rect 98992 25540 99016 25542
rect 99072 25540 99096 25542
rect 99152 25540 99176 25542
rect 99232 25540 99238 25542
rect 98930 25531 99238 25540
rect 99288 25356 99340 25362
rect 99288 25298 99340 25304
rect 98930 24508 99238 24517
rect 98930 24506 98936 24508
rect 98992 24506 99016 24508
rect 99072 24506 99096 24508
rect 99152 24506 99176 24508
rect 99232 24506 99238 24508
rect 98992 24454 98994 24506
rect 99174 24454 99176 24506
rect 98930 24452 98936 24454
rect 98992 24452 99016 24454
rect 99072 24452 99096 24454
rect 99152 24452 99176 24454
rect 99232 24452 99238 24454
rect 98930 24443 99238 24452
rect 99300 23866 99328 25298
rect 99380 24744 99432 24750
rect 99380 24686 99432 24692
rect 99288 23860 99340 23866
rect 99288 23802 99340 23808
rect 98930 23420 99238 23429
rect 98930 23418 98936 23420
rect 98992 23418 99016 23420
rect 99072 23418 99096 23420
rect 99152 23418 99176 23420
rect 99232 23418 99238 23420
rect 98992 23366 98994 23418
rect 99174 23366 99176 23418
rect 98930 23364 98936 23366
rect 98992 23364 99016 23366
rect 99072 23364 99096 23366
rect 99152 23364 99176 23366
rect 99232 23364 99238 23366
rect 98930 23355 99238 23364
rect 99392 22778 99420 24686
rect 99472 23724 99524 23730
rect 99472 23666 99524 23672
rect 99484 22778 99512 23666
rect 99380 22772 99432 22778
rect 99380 22714 99432 22720
rect 99472 22772 99524 22778
rect 99472 22714 99524 22720
rect 99288 22636 99340 22642
rect 99288 22578 99340 22584
rect 98828 22432 98880 22438
rect 98828 22374 98880 22380
rect 98930 22332 99238 22341
rect 98930 22330 98936 22332
rect 98992 22330 99016 22332
rect 99072 22330 99096 22332
rect 99152 22330 99176 22332
rect 99232 22330 99238 22332
rect 98992 22278 98994 22330
rect 99174 22278 99176 22330
rect 98930 22276 98936 22278
rect 98992 22276 99016 22278
rect 99072 22276 99096 22278
rect 99152 22276 99176 22278
rect 99232 22276 99238 22278
rect 98930 22267 99238 22276
rect 98736 21956 98788 21962
rect 98736 21898 98788 21904
rect 99300 21894 99328 22578
rect 99380 22432 99432 22438
rect 99380 22374 99432 22380
rect 98644 21888 98696 21894
rect 98644 21830 98696 21836
rect 99288 21888 99340 21894
rect 99288 21830 99340 21836
rect 98656 18222 98684 21830
rect 98930 21244 99238 21253
rect 98930 21242 98936 21244
rect 98992 21242 99016 21244
rect 99072 21242 99096 21244
rect 99152 21242 99176 21244
rect 99232 21242 99238 21244
rect 98992 21190 98994 21242
rect 99174 21190 99176 21242
rect 98930 21188 98936 21190
rect 98992 21188 99016 21190
rect 99072 21188 99096 21190
rect 99152 21188 99176 21190
rect 99232 21188 99238 21190
rect 98930 21179 99238 21188
rect 98930 20156 99238 20165
rect 98930 20154 98936 20156
rect 98992 20154 99016 20156
rect 99072 20154 99096 20156
rect 99152 20154 99176 20156
rect 99232 20154 99238 20156
rect 98992 20102 98994 20154
rect 99174 20102 99176 20154
rect 98930 20100 98936 20102
rect 98992 20100 99016 20102
rect 99072 20100 99096 20102
rect 99152 20100 99176 20102
rect 99232 20100 99238 20102
rect 98930 20091 99238 20100
rect 98828 19916 98880 19922
rect 98828 19858 98880 19864
rect 98840 18222 98868 19858
rect 98930 19068 99238 19077
rect 98930 19066 98936 19068
rect 98992 19066 99016 19068
rect 99072 19066 99096 19068
rect 99152 19066 99176 19068
rect 99232 19066 99238 19068
rect 98992 19014 98994 19066
rect 99174 19014 99176 19066
rect 98930 19012 98936 19014
rect 98992 19012 99016 19014
rect 99072 19012 99096 19014
rect 99152 19012 99176 19014
rect 99232 19012 99238 19014
rect 98930 19003 99238 19012
rect 98644 18216 98696 18222
rect 98644 18158 98696 18164
rect 98828 18216 98880 18222
rect 98828 18158 98880 18164
rect 98930 17980 99238 17989
rect 98930 17978 98936 17980
rect 98992 17978 99016 17980
rect 99072 17978 99096 17980
rect 99152 17978 99176 17980
rect 99232 17978 99238 17980
rect 98992 17926 98994 17978
rect 99174 17926 99176 17978
rect 98930 17924 98936 17926
rect 98992 17924 99016 17926
rect 99072 17924 99096 17926
rect 99152 17924 99176 17926
rect 99232 17924 99238 17926
rect 98930 17915 99238 17924
rect 99392 17377 99420 22374
rect 99484 22234 99512 22714
rect 99576 22438 99604 25842
rect 99666 25052 99974 25061
rect 99666 25050 99672 25052
rect 99728 25050 99752 25052
rect 99808 25050 99832 25052
rect 99888 25050 99912 25052
rect 99968 25050 99974 25052
rect 99728 24998 99730 25050
rect 99910 24998 99912 25050
rect 99666 24996 99672 24998
rect 99728 24996 99752 24998
rect 99808 24996 99832 24998
rect 99888 24996 99912 24998
rect 99968 24996 99974 24998
rect 99666 24987 99974 24996
rect 99666 23964 99974 23973
rect 99666 23962 99672 23964
rect 99728 23962 99752 23964
rect 99808 23962 99832 23964
rect 99888 23962 99912 23964
rect 99968 23962 99974 23964
rect 99728 23910 99730 23962
rect 99910 23910 99912 23962
rect 99666 23908 99672 23910
rect 99728 23908 99752 23910
rect 99808 23908 99832 23910
rect 99888 23908 99912 23910
rect 99968 23908 99974 23910
rect 99666 23899 99974 23908
rect 100036 23730 100064 25978
rect 100220 25294 100248 30670
rect 100312 29102 100340 35866
rect 100300 29096 100352 29102
rect 100300 29038 100352 29044
rect 100312 27470 100340 29038
rect 100300 27464 100352 27470
rect 100300 27406 100352 27412
rect 100484 26376 100536 26382
rect 100484 26318 100536 26324
rect 100496 25945 100524 26318
rect 100482 25936 100538 25945
rect 100482 25871 100538 25880
rect 100208 25288 100260 25294
rect 100208 25230 100260 25236
rect 100220 24750 100248 25230
rect 100208 24744 100260 24750
rect 100208 24686 100260 24692
rect 100024 23724 100076 23730
rect 100024 23666 100076 23672
rect 99666 22876 99974 22885
rect 99666 22874 99672 22876
rect 99728 22874 99752 22876
rect 99808 22874 99832 22876
rect 99888 22874 99912 22876
rect 99968 22874 99974 22876
rect 99728 22822 99730 22874
rect 99910 22822 99912 22874
rect 99666 22820 99672 22822
rect 99728 22820 99752 22822
rect 99808 22820 99832 22822
rect 99888 22820 99912 22822
rect 99968 22820 99974 22822
rect 99666 22811 99974 22820
rect 99564 22432 99616 22438
rect 99564 22374 99616 22380
rect 99472 22228 99524 22234
rect 99472 22170 99524 22176
rect 99666 21788 99974 21797
rect 99666 21786 99672 21788
rect 99728 21786 99752 21788
rect 99808 21786 99832 21788
rect 99888 21786 99912 21788
rect 99968 21786 99974 21788
rect 99728 21734 99730 21786
rect 99910 21734 99912 21786
rect 99666 21732 99672 21734
rect 99728 21732 99752 21734
rect 99808 21732 99832 21734
rect 99888 21732 99912 21734
rect 99968 21732 99974 21734
rect 99666 21723 99974 21732
rect 99666 20700 99974 20709
rect 99666 20698 99672 20700
rect 99728 20698 99752 20700
rect 99808 20698 99832 20700
rect 99888 20698 99912 20700
rect 99968 20698 99974 20700
rect 99728 20646 99730 20698
rect 99910 20646 99912 20698
rect 99666 20644 99672 20646
rect 99728 20644 99752 20646
rect 99808 20644 99832 20646
rect 99888 20644 99912 20646
rect 99968 20644 99974 20646
rect 99666 20635 99974 20644
rect 100220 19922 100248 24686
rect 100208 19916 100260 19922
rect 100208 19858 100260 19864
rect 99666 19612 99974 19621
rect 99666 19610 99672 19612
rect 99728 19610 99752 19612
rect 99808 19610 99832 19612
rect 99888 19610 99912 19612
rect 99968 19610 99974 19612
rect 99728 19558 99730 19610
rect 99910 19558 99912 19610
rect 99666 19556 99672 19558
rect 99728 19556 99752 19558
rect 99808 19556 99832 19558
rect 99888 19556 99912 19558
rect 99968 19556 99974 19558
rect 99666 19547 99974 19556
rect 99666 18524 99974 18533
rect 99666 18522 99672 18524
rect 99728 18522 99752 18524
rect 99808 18522 99832 18524
rect 99888 18522 99912 18524
rect 99968 18522 99974 18524
rect 99728 18470 99730 18522
rect 99910 18470 99912 18522
rect 99666 18468 99672 18470
rect 99728 18468 99752 18470
rect 99808 18468 99832 18470
rect 99888 18468 99912 18470
rect 99968 18468 99974 18470
rect 99666 18459 99974 18468
rect 99666 17436 99974 17445
rect 99666 17434 99672 17436
rect 99728 17434 99752 17436
rect 99808 17434 99832 17436
rect 99888 17434 99912 17436
rect 99968 17434 99974 17436
rect 99728 17382 99730 17434
rect 99910 17382 99912 17434
rect 99666 17380 99672 17382
rect 99728 17380 99752 17382
rect 99808 17380 99832 17382
rect 99888 17380 99912 17382
rect 99968 17380 99974 17382
rect 99378 17368 99434 17377
rect 99666 17371 99974 17380
rect 99378 17303 99434 17312
rect 98930 16892 99238 16901
rect 98930 16890 98936 16892
rect 98992 16890 99016 16892
rect 99072 16890 99096 16892
rect 99152 16890 99176 16892
rect 99232 16890 99238 16892
rect 98992 16838 98994 16890
rect 99174 16838 99176 16890
rect 98930 16836 98936 16838
rect 98992 16836 99016 16838
rect 99072 16836 99096 16838
rect 99152 16836 99176 16838
rect 99232 16836 99238 16838
rect 98930 16827 99238 16836
rect 99666 16348 99974 16357
rect 99666 16346 99672 16348
rect 99728 16346 99752 16348
rect 99808 16346 99832 16348
rect 99888 16346 99912 16348
rect 99968 16346 99974 16348
rect 99728 16294 99730 16346
rect 99910 16294 99912 16346
rect 99666 16292 99672 16294
rect 99728 16292 99752 16294
rect 99808 16292 99832 16294
rect 99888 16292 99912 16294
rect 99968 16292 99974 16294
rect 98550 16280 98606 16289
rect 99666 16283 99974 16292
rect 98550 16215 98606 16224
rect 98930 15804 99238 15813
rect 98930 15802 98936 15804
rect 98992 15802 99016 15804
rect 99072 15802 99096 15804
rect 99152 15802 99176 15804
rect 99232 15802 99238 15804
rect 98992 15750 98994 15802
rect 99174 15750 99176 15802
rect 98930 15748 98936 15750
rect 98992 15748 99016 15750
rect 99072 15748 99096 15750
rect 99152 15748 99176 15750
rect 99232 15748 99238 15750
rect 98930 15739 99238 15748
rect 99666 15260 99974 15269
rect 99666 15258 99672 15260
rect 99728 15258 99752 15260
rect 99808 15258 99832 15260
rect 99888 15258 99912 15260
rect 99968 15258 99974 15260
rect 99728 15206 99730 15258
rect 99910 15206 99912 15258
rect 99666 15204 99672 15206
rect 99728 15204 99752 15206
rect 99808 15204 99832 15206
rect 99888 15204 99912 15206
rect 99968 15204 99974 15206
rect 99666 15195 99974 15204
rect 98930 14716 99238 14725
rect 98930 14714 98936 14716
rect 98992 14714 99016 14716
rect 99072 14714 99096 14716
rect 99152 14714 99176 14716
rect 99232 14714 99238 14716
rect 98992 14662 98994 14714
rect 99174 14662 99176 14714
rect 98930 14660 98936 14662
rect 98992 14660 99016 14662
rect 99072 14660 99096 14662
rect 99152 14660 99176 14662
rect 99232 14660 99238 14662
rect 98930 14651 99238 14660
rect 99666 14172 99974 14181
rect 99666 14170 99672 14172
rect 99728 14170 99752 14172
rect 99808 14170 99832 14172
rect 99888 14170 99912 14172
rect 99968 14170 99974 14172
rect 99728 14118 99730 14170
rect 99910 14118 99912 14170
rect 99666 14116 99672 14118
rect 99728 14116 99752 14118
rect 99808 14116 99832 14118
rect 99888 14116 99912 14118
rect 99968 14116 99974 14118
rect 99666 14107 99974 14116
rect 98930 13628 99238 13637
rect 98930 13626 98936 13628
rect 98992 13626 99016 13628
rect 99072 13626 99096 13628
rect 99152 13626 99176 13628
rect 99232 13626 99238 13628
rect 98992 13574 98994 13626
rect 99174 13574 99176 13626
rect 98930 13572 98936 13574
rect 98992 13572 99016 13574
rect 99072 13572 99096 13574
rect 99152 13572 99176 13574
rect 99232 13572 99238 13574
rect 98930 13563 99238 13572
rect 99666 13084 99974 13093
rect 99666 13082 99672 13084
rect 99728 13082 99752 13084
rect 99808 13082 99832 13084
rect 99888 13082 99912 13084
rect 99968 13082 99974 13084
rect 99728 13030 99730 13082
rect 99910 13030 99912 13082
rect 99666 13028 99672 13030
rect 99728 13028 99752 13030
rect 99808 13028 99832 13030
rect 99888 13028 99912 13030
rect 99968 13028 99974 13030
rect 99666 13019 99974 13028
rect 98930 12540 99238 12549
rect 98930 12538 98936 12540
rect 98992 12538 99016 12540
rect 99072 12538 99096 12540
rect 99152 12538 99176 12540
rect 99232 12538 99238 12540
rect 98992 12486 98994 12538
rect 99174 12486 99176 12538
rect 98930 12484 98936 12486
rect 98992 12484 99016 12486
rect 99072 12484 99096 12486
rect 99152 12484 99176 12486
rect 99232 12484 99238 12486
rect 98930 12475 99238 12484
rect 99666 11996 99974 12005
rect 99666 11994 99672 11996
rect 99728 11994 99752 11996
rect 99808 11994 99832 11996
rect 99888 11994 99912 11996
rect 99968 11994 99974 11996
rect 99728 11942 99730 11994
rect 99910 11942 99912 11994
rect 99666 11940 99672 11942
rect 99728 11940 99752 11942
rect 99808 11940 99832 11942
rect 99888 11940 99912 11942
rect 99968 11940 99974 11942
rect 99666 11931 99974 11940
rect 98930 11452 99238 11461
rect 98930 11450 98936 11452
rect 98992 11450 99016 11452
rect 99072 11450 99096 11452
rect 99152 11450 99176 11452
rect 99232 11450 99238 11452
rect 98992 11398 98994 11450
rect 99174 11398 99176 11450
rect 98930 11396 98936 11398
rect 98992 11396 99016 11398
rect 99072 11396 99096 11398
rect 99152 11396 99176 11398
rect 99232 11396 99238 11398
rect 98930 11387 99238 11396
rect 99666 10908 99974 10917
rect 99666 10906 99672 10908
rect 99728 10906 99752 10908
rect 99808 10906 99832 10908
rect 99888 10906 99912 10908
rect 99968 10906 99974 10908
rect 99728 10854 99730 10906
rect 99910 10854 99912 10906
rect 99666 10852 99672 10854
rect 99728 10852 99752 10854
rect 99808 10852 99832 10854
rect 99888 10852 99912 10854
rect 99968 10852 99974 10854
rect 99666 10843 99974 10852
rect 98930 10364 99238 10373
rect 98930 10362 98936 10364
rect 98992 10362 99016 10364
rect 99072 10362 99096 10364
rect 99152 10362 99176 10364
rect 99232 10362 99238 10364
rect 98992 10310 98994 10362
rect 99174 10310 99176 10362
rect 98930 10308 98936 10310
rect 98992 10308 99016 10310
rect 99072 10308 99096 10310
rect 99152 10308 99176 10310
rect 99232 10308 99238 10310
rect 98930 10299 99238 10308
rect 99666 9820 99974 9829
rect 99666 9818 99672 9820
rect 99728 9818 99752 9820
rect 99808 9818 99832 9820
rect 99888 9818 99912 9820
rect 99968 9818 99974 9820
rect 99728 9766 99730 9818
rect 99910 9766 99912 9818
rect 99666 9764 99672 9766
rect 99728 9764 99752 9766
rect 99808 9764 99832 9766
rect 99888 9764 99912 9766
rect 99968 9764 99974 9766
rect 99666 9755 99974 9764
rect 98930 9276 99238 9285
rect 98930 9274 98936 9276
rect 98992 9274 99016 9276
rect 99072 9274 99096 9276
rect 99152 9274 99176 9276
rect 99232 9274 99238 9276
rect 98992 9222 98994 9274
rect 99174 9222 99176 9274
rect 98930 9220 98936 9222
rect 98992 9220 99016 9222
rect 99072 9220 99096 9222
rect 99152 9220 99176 9222
rect 99232 9220 99238 9222
rect 98930 9211 99238 9220
rect 99666 8732 99974 8741
rect 99666 8730 99672 8732
rect 99728 8730 99752 8732
rect 99808 8730 99832 8732
rect 99888 8730 99912 8732
rect 99968 8730 99974 8732
rect 99728 8678 99730 8730
rect 99910 8678 99912 8730
rect 99666 8676 99672 8678
rect 99728 8676 99752 8678
rect 99808 8676 99832 8678
rect 99888 8676 99912 8678
rect 99968 8676 99974 8678
rect 99666 8667 99974 8676
rect 98930 8188 99238 8197
rect 98930 8186 98936 8188
rect 98992 8186 99016 8188
rect 99072 8186 99096 8188
rect 99152 8186 99176 8188
rect 99232 8186 99238 8188
rect 98992 8134 98994 8186
rect 99174 8134 99176 8186
rect 98930 8132 98936 8134
rect 98992 8132 99016 8134
rect 99072 8132 99096 8134
rect 99152 8132 99176 8134
rect 99232 8132 99238 8134
rect 98930 8123 99238 8132
rect 99666 7644 99974 7653
rect 99666 7642 99672 7644
rect 99728 7642 99752 7644
rect 99808 7642 99832 7644
rect 99888 7642 99912 7644
rect 99968 7642 99974 7644
rect 99728 7590 99730 7642
rect 99910 7590 99912 7642
rect 99666 7588 99672 7590
rect 99728 7588 99752 7590
rect 99808 7588 99832 7590
rect 99888 7588 99912 7590
rect 99968 7588 99974 7590
rect 99666 7579 99974 7588
rect 98930 7100 99238 7109
rect 98930 7098 98936 7100
rect 98992 7098 99016 7100
rect 99072 7098 99096 7100
rect 99152 7098 99176 7100
rect 99232 7098 99238 7100
rect 98992 7046 98994 7098
rect 99174 7046 99176 7098
rect 98930 7044 98936 7046
rect 98992 7044 99016 7046
rect 99072 7044 99096 7046
rect 99152 7044 99176 7046
rect 99232 7044 99238 7046
rect 98930 7035 99238 7044
rect 98012 6886 98408 6914
rect 98012 3913 98040 6886
rect 99666 6556 99974 6565
rect 99666 6554 99672 6556
rect 99728 6554 99752 6556
rect 99808 6554 99832 6556
rect 99888 6554 99912 6556
rect 99968 6554 99974 6556
rect 99728 6502 99730 6554
rect 99910 6502 99912 6554
rect 99666 6500 99672 6502
rect 99728 6500 99752 6502
rect 99808 6500 99832 6502
rect 99888 6500 99912 6502
rect 99968 6500 99974 6502
rect 99666 6491 99974 6500
rect 98930 6012 99238 6021
rect 98930 6010 98936 6012
rect 98992 6010 99016 6012
rect 99072 6010 99096 6012
rect 99152 6010 99176 6012
rect 99232 6010 99238 6012
rect 98992 5958 98994 6010
rect 99174 5958 99176 6010
rect 98930 5956 98936 5958
rect 98992 5956 99016 5958
rect 99072 5956 99096 5958
rect 99152 5956 99176 5958
rect 99232 5956 99238 5958
rect 98930 5947 99238 5956
rect 99666 5468 99974 5477
rect 99666 5466 99672 5468
rect 99728 5466 99752 5468
rect 99808 5466 99832 5468
rect 99888 5466 99912 5468
rect 99968 5466 99974 5468
rect 99728 5414 99730 5466
rect 99910 5414 99912 5466
rect 99666 5412 99672 5414
rect 99728 5412 99752 5414
rect 99808 5412 99832 5414
rect 99888 5412 99912 5414
rect 99968 5412 99974 5414
rect 99666 5403 99974 5412
rect 98930 4924 99238 4933
rect 98930 4922 98936 4924
rect 98992 4922 99016 4924
rect 99072 4922 99096 4924
rect 99152 4922 99176 4924
rect 99232 4922 99238 4924
rect 98992 4870 98994 4922
rect 99174 4870 99176 4922
rect 98930 4868 98936 4870
rect 98992 4868 99016 4870
rect 99072 4868 99096 4870
rect 99152 4868 99176 4870
rect 99232 4868 99238 4870
rect 98930 4859 99238 4868
rect 99666 4380 99974 4389
rect 99666 4378 99672 4380
rect 99728 4378 99752 4380
rect 99808 4378 99832 4380
rect 99888 4378 99912 4380
rect 99968 4378 99974 4380
rect 99728 4326 99730 4378
rect 99910 4326 99912 4378
rect 99666 4324 99672 4326
rect 99728 4324 99752 4326
rect 99808 4324 99832 4326
rect 99888 4324 99912 4326
rect 99968 4324 99974 4326
rect 99666 4315 99974 4324
rect 97998 3904 98054 3913
rect 97998 3839 98054 3848
rect 98930 3836 99238 3845
rect 98930 3834 98936 3836
rect 98992 3834 99016 3836
rect 99072 3834 99096 3836
rect 99152 3834 99176 3836
rect 99232 3834 99238 3836
rect 98992 3782 98994 3834
rect 99174 3782 99176 3834
rect 98930 3780 98936 3782
rect 98992 3780 99016 3782
rect 99072 3780 99096 3782
rect 99152 3780 99176 3782
rect 99232 3780 99238 3782
rect 97538 3768 97594 3777
rect 98930 3771 99238 3780
rect 97538 3703 97594 3712
rect 97354 3632 97410 3641
rect 97354 3567 97410 3576
rect 17406 3496 17462 3505
rect 17406 3431 17462 3440
rect 19982 3496 20038 3505
rect 19982 3431 20038 3440
rect 20626 3496 20682 3505
rect 20626 3431 20682 3440
rect 21914 3496 21970 3505
rect 21914 3431 21970 3440
rect 24490 3496 24546 3505
rect 24490 3431 24546 3440
rect 25778 3496 25834 3505
rect 25778 3431 25834 3440
rect 27066 3496 27122 3505
rect 27066 3431 27122 3440
rect 27710 3496 27766 3505
rect 27710 3431 27766 3440
rect 30286 3496 30342 3505
rect 30286 3431 30342 3440
rect 33506 3496 33562 3505
rect 33506 3431 33562 3440
rect 34794 3496 34850 3505
rect 34794 3431 34850 3440
rect 1680 3292 1816 3301
rect 1736 3290 1760 3292
rect 1742 3238 1754 3290
rect 1736 3236 1760 3238
rect 1680 3227 1816 3236
rect 1312 2748 1448 2757
rect 1368 2746 1392 2748
rect 1374 2694 1386 2746
rect 1368 2692 1392 2694
rect 1312 2683 1448 2692
rect 1680 2204 1816 2213
rect 1736 2202 1760 2204
rect 1742 2150 1754 2202
rect 1736 2148 1760 2150
rect 1680 2139 1816 2148
rect 17420 800 17448 3431
rect 18694 2816 18750 2825
rect 18694 2751 18750 2760
rect 18708 800 18736 2751
rect 19996 800 20024 3431
rect 20640 800 20668 3431
rect 21928 800 21956 3431
rect 23202 2816 23258 2825
rect 23202 2751 23258 2760
rect 23216 800 23244 2751
rect 24504 800 24532 3431
rect 25792 800 25820 3431
rect 27080 800 27108 3431
rect 27724 800 27752 3431
rect 28998 2816 29054 2825
rect 28998 2751 29054 2760
rect 29012 800 29040 2751
rect 30300 800 30328 3431
rect 31574 2816 31630 2825
rect 31574 2751 31630 2760
rect 32862 2816 32918 2825
rect 32862 2751 32918 2760
rect 31588 800 31616 2751
rect 32876 800 32904 2751
rect 33520 800 33548 3431
rect 34808 800 34836 3431
rect 99666 3292 99974 3301
rect 99666 3290 99672 3292
rect 99728 3290 99752 3292
rect 99808 3290 99832 3292
rect 99888 3290 99912 3292
rect 99968 3290 99974 3292
rect 99728 3238 99730 3290
rect 99910 3238 99912 3290
rect 99666 3236 99672 3238
rect 99728 3236 99752 3238
rect 99808 3236 99832 3238
rect 99888 3236 99912 3238
rect 99968 3236 99974 3238
rect 99666 3227 99974 3236
rect 36082 2816 36138 2825
rect 36082 2751 36138 2760
rect 37370 2816 37426 2825
rect 37370 2751 37426 2760
rect 36096 800 36124 2751
rect 37384 800 37412 2751
rect 98930 2748 99238 2757
rect 98930 2746 98936 2748
rect 98992 2746 99016 2748
rect 99072 2746 99096 2748
rect 99152 2746 99176 2748
rect 99232 2746 99238 2748
rect 98992 2694 98994 2746
rect 99174 2694 99176 2746
rect 98930 2692 98936 2694
rect 98992 2692 99016 2694
rect 99072 2692 99096 2694
rect 99152 2692 99176 2694
rect 99232 2692 99238 2694
rect 98930 2683 99238 2692
rect 99666 2204 99974 2213
rect 99666 2202 99672 2204
rect 99728 2202 99752 2204
rect 99808 2202 99832 2204
rect 99888 2202 99912 2204
rect 99968 2202 99974 2204
rect 99728 2150 99730 2202
rect 99910 2150 99912 2202
rect 99666 2148 99672 2150
rect 99728 2148 99752 2150
rect 99808 2148 99832 2150
rect 99888 2148 99912 2150
rect 99968 2148 99974 2150
rect 99666 2139 99974 2148
rect 17406 0 17462 800
rect 18694 0 18750 800
rect 19982 0 20038 800
rect 20626 0 20682 800
rect 21914 0 21970 800
rect 23202 0 23258 800
rect 24490 0 24546 800
rect 25778 0 25834 800
rect 27066 0 27122 800
rect 27710 0 27766 800
rect 28998 0 29054 800
rect 30286 0 30342 800
rect 31574 0 31630 800
rect 32862 0 32918 800
rect 33506 0 33562 800
rect 34794 0 34850 800
rect 36082 0 36138 800
rect 37370 0 37426 800
<< via2 >>
rect 4220 101754 4276 101756
rect 4300 101754 4356 101756
rect 4380 101754 4436 101756
rect 4460 101754 4516 101756
rect 4220 101702 4266 101754
rect 4266 101702 4276 101754
rect 4300 101702 4330 101754
rect 4330 101702 4342 101754
rect 4342 101702 4356 101754
rect 4380 101702 4394 101754
rect 4394 101702 4406 101754
rect 4406 101702 4436 101754
rect 4460 101702 4470 101754
rect 4470 101702 4516 101754
rect 4220 101700 4276 101702
rect 4300 101700 4356 101702
rect 4380 101700 4436 101702
rect 4460 101700 4516 101702
rect 34940 101754 34996 101756
rect 35020 101754 35076 101756
rect 35100 101754 35156 101756
rect 35180 101754 35236 101756
rect 34940 101702 34986 101754
rect 34986 101702 34996 101754
rect 35020 101702 35050 101754
rect 35050 101702 35062 101754
rect 35062 101702 35076 101754
rect 35100 101702 35114 101754
rect 35114 101702 35126 101754
rect 35126 101702 35156 101754
rect 35180 101702 35190 101754
rect 35190 101702 35236 101754
rect 34940 101700 34996 101702
rect 35020 101700 35076 101702
rect 35100 101700 35156 101702
rect 35180 101700 35236 101702
rect 65660 101754 65716 101756
rect 65740 101754 65796 101756
rect 65820 101754 65876 101756
rect 65900 101754 65956 101756
rect 65660 101702 65706 101754
rect 65706 101702 65716 101754
rect 65740 101702 65770 101754
rect 65770 101702 65782 101754
rect 65782 101702 65796 101754
rect 65820 101702 65834 101754
rect 65834 101702 65846 101754
rect 65846 101702 65876 101754
rect 65900 101702 65910 101754
rect 65910 101702 65956 101754
rect 65660 101700 65716 101702
rect 65740 101700 65796 101702
rect 65820 101700 65876 101702
rect 65900 101700 65956 101702
rect 96380 101754 96436 101756
rect 96460 101754 96516 101756
rect 96540 101754 96596 101756
rect 96620 101754 96676 101756
rect 96380 101702 96426 101754
rect 96426 101702 96436 101754
rect 96460 101702 96490 101754
rect 96490 101702 96502 101754
rect 96502 101702 96516 101754
rect 96540 101702 96554 101754
rect 96554 101702 96566 101754
rect 96566 101702 96596 101754
rect 96620 101702 96630 101754
rect 96630 101702 96676 101754
rect 96380 101700 96436 101702
rect 96460 101700 96516 101702
rect 96540 101700 96596 101702
rect 96620 101700 96676 101702
rect 4880 101210 4936 101212
rect 4960 101210 5016 101212
rect 5040 101210 5096 101212
rect 5120 101210 5176 101212
rect 4880 101158 4926 101210
rect 4926 101158 4936 101210
rect 4960 101158 4990 101210
rect 4990 101158 5002 101210
rect 5002 101158 5016 101210
rect 5040 101158 5054 101210
rect 5054 101158 5066 101210
rect 5066 101158 5096 101210
rect 5120 101158 5130 101210
rect 5130 101158 5176 101210
rect 4880 101156 4936 101158
rect 4960 101156 5016 101158
rect 5040 101156 5096 101158
rect 5120 101156 5176 101158
rect 35600 101210 35656 101212
rect 35680 101210 35736 101212
rect 35760 101210 35816 101212
rect 35840 101210 35896 101212
rect 35600 101158 35646 101210
rect 35646 101158 35656 101210
rect 35680 101158 35710 101210
rect 35710 101158 35722 101210
rect 35722 101158 35736 101210
rect 35760 101158 35774 101210
rect 35774 101158 35786 101210
rect 35786 101158 35816 101210
rect 35840 101158 35850 101210
rect 35850 101158 35896 101210
rect 35600 101156 35656 101158
rect 35680 101156 35736 101158
rect 35760 101156 35816 101158
rect 35840 101156 35896 101158
rect 4220 100666 4276 100668
rect 4300 100666 4356 100668
rect 4380 100666 4436 100668
rect 4460 100666 4516 100668
rect 4220 100614 4266 100666
rect 4266 100614 4276 100666
rect 4300 100614 4330 100666
rect 4330 100614 4342 100666
rect 4342 100614 4356 100666
rect 4380 100614 4394 100666
rect 4394 100614 4406 100666
rect 4406 100614 4436 100666
rect 4460 100614 4470 100666
rect 4470 100614 4516 100666
rect 4220 100612 4276 100614
rect 4300 100612 4356 100614
rect 4380 100612 4436 100614
rect 4460 100612 4516 100614
rect 34940 100666 34996 100668
rect 35020 100666 35076 100668
rect 35100 100666 35156 100668
rect 35180 100666 35236 100668
rect 34940 100614 34986 100666
rect 34986 100614 34996 100666
rect 35020 100614 35050 100666
rect 35050 100614 35062 100666
rect 35062 100614 35076 100666
rect 35100 100614 35114 100666
rect 35114 100614 35126 100666
rect 35126 100614 35156 100666
rect 35180 100614 35190 100666
rect 35190 100614 35236 100666
rect 34940 100612 34996 100614
rect 35020 100612 35076 100614
rect 35100 100612 35156 100614
rect 35180 100612 35236 100614
rect 4880 100122 4936 100124
rect 4960 100122 5016 100124
rect 5040 100122 5096 100124
rect 5120 100122 5176 100124
rect 4880 100070 4926 100122
rect 4926 100070 4936 100122
rect 4960 100070 4990 100122
rect 4990 100070 5002 100122
rect 5002 100070 5016 100122
rect 5040 100070 5054 100122
rect 5054 100070 5066 100122
rect 5066 100070 5096 100122
rect 5120 100070 5130 100122
rect 5130 100070 5176 100122
rect 4880 100068 4936 100070
rect 4960 100068 5016 100070
rect 5040 100068 5096 100070
rect 5120 100068 5176 100070
rect 35600 100122 35656 100124
rect 35680 100122 35736 100124
rect 35760 100122 35816 100124
rect 35840 100122 35896 100124
rect 35600 100070 35646 100122
rect 35646 100070 35656 100122
rect 35680 100070 35710 100122
rect 35710 100070 35722 100122
rect 35722 100070 35736 100122
rect 35760 100070 35774 100122
rect 35774 100070 35786 100122
rect 35786 100070 35816 100122
rect 35840 100070 35850 100122
rect 35850 100070 35896 100122
rect 35600 100068 35656 100070
rect 35680 100068 35736 100070
rect 35760 100068 35816 100070
rect 35840 100068 35896 100070
rect 4220 99578 4276 99580
rect 4300 99578 4356 99580
rect 4380 99578 4436 99580
rect 4460 99578 4516 99580
rect 4220 99526 4266 99578
rect 4266 99526 4276 99578
rect 4300 99526 4330 99578
rect 4330 99526 4342 99578
rect 4342 99526 4356 99578
rect 4380 99526 4394 99578
rect 4394 99526 4406 99578
rect 4406 99526 4436 99578
rect 4460 99526 4470 99578
rect 4470 99526 4516 99578
rect 4220 99524 4276 99526
rect 4300 99524 4356 99526
rect 4380 99524 4436 99526
rect 4460 99524 4516 99526
rect 34940 99578 34996 99580
rect 35020 99578 35076 99580
rect 35100 99578 35156 99580
rect 35180 99578 35236 99580
rect 34940 99526 34986 99578
rect 34986 99526 34996 99578
rect 35020 99526 35050 99578
rect 35050 99526 35062 99578
rect 35062 99526 35076 99578
rect 35100 99526 35114 99578
rect 35114 99526 35126 99578
rect 35126 99526 35156 99578
rect 35180 99526 35190 99578
rect 35190 99526 35236 99578
rect 34940 99524 34996 99526
rect 35020 99524 35076 99526
rect 35100 99524 35156 99526
rect 35180 99524 35236 99526
rect 4880 99034 4936 99036
rect 4960 99034 5016 99036
rect 5040 99034 5096 99036
rect 5120 99034 5176 99036
rect 4880 98982 4926 99034
rect 4926 98982 4936 99034
rect 4960 98982 4990 99034
rect 4990 98982 5002 99034
rect 5002 98982 5016 99034
rect 5040 98982 5054 99034
rect 5054 98982 5066 99034
rect 5066 98982 5096 99034
rect 5120 98982 5130 99034
rect 5130 98982 5176 99034
rect 4880 98980 4936 98982
rect 4960 98980 5016 98982
rect 5040 98980 5096 98982
rect 5120 98980 5176 98982
rect 35600 99034 35656 99036
rect 35680 99034 35736 99036
rect 35760 99034 35816 99036
rect 35840 99034 35896 99036
rect 35600 98982 35646 99034
rect 35646 98982 35656 99034
rect 35680 98982 35710 99034
rect 35710 98982 35722 99034
rect 35722 98982 35736 99034
rect 35760 98982 35774 99034
rect 35774 98982 35786 99034
rect 35786 98982 35816 99034
rect 35840 98982 35850 99034
rect 35850 98982 35896 99034
rect 35600 98980 35656 98982
rect 35680 98980 35736 98982
rect 35760 98980 35816 98982
rect 35840 98980 35896 98982
rect 4220 98490 4276 98492
rect 4300 98490 4356 98492
rect 4380 98490 4436 98492
rect 4460 98490 4516 98492
rect 4220 98438 4266 98490
rect 4266 98438 4276 98490
rect 4300 98438 4330 98490
rect 4330 98438 4342 98490
rect 4342 98438 4356 98490
rect 4380 98438 4394 98490
rect 4394 98438 4406 98490
rect 4406 98438 4436 98490
rect 4460 98438 4470 98490
rect 4470 98438 4516 98490
rect 4220 98436 4276 98438
rect 4300 98436 4356 98438
rect 4380 98436 4436 98438
rect 4460 98436 4516 98438
rect 34940 98490 34996 98492
rect 35020 98490 35076 98492
rect 35100 98490 35156 98492
rect 35180 98490 35236 98492
rect 34940 98438 34986 98490
rect 34986 98438 34996 98490
rect 35020 98438 35050 98490
rect 35050 98438 35062 98490
rect 35062 98438 35076 98490
rect 35100 98438 35114 98490
rect 35114 98438 35126 98490
rect 35126 98438 35156 98490
rect 35180 98438 35190 98490
rect 35190 98438 35236 98490
rect 34940 98436 34996 98438
rect 35020 98436 35076 98438
rect 35100 98436 35156 98438
rect 35180 98436 35236 98438
rect 4880 97946 4936 97948
rect 4960 97946 5016 97948
rect 5040 97946 5096 97948
rect 5120 97946 5176 97948
rect 4880 97894 4926 97946
rect 4926 97894 4936 97946
rect 4960 97894 4990 97946
rect 4990 97894 5002 97946
rect 5002 97894 5016 97946
rect 5040 97894 5054 97946
rect 5054 97894 5066 97946
rect 5066 97894 5096 97946
rect 5120 97894 5130 97946
rect 5130 97894 5176 97946
rect 4880 97892 4936 97894
rect 4960 97892 5016 97894
rect 5040 97892 5096 97894
rect 5120 97892 5176 97894
rect 35600 97946 35656 97948
rect 35680 97946 35736 97948
rect 35760 97946 35816 97948
rect 35840 97946 35896 97948
rect 35600 97894 35646 97946
rect 35646 97894 35656 97946
rect 35680 97894 35710 97946
rect 35710 97894 35722 97946
rect 35722 97894 35736 97946
rect 35760 97894 35774 97946
rect 35774 97894 35786 97946
rect 35786 97894 35816 97946
rect 35840 97894 35850 97946
rect 35850 97894 35896 97946
rect 35600 97892 35656 97894
rect 35680 97892 35736 97894
rect 35760 97892 35816 97894
rect 35840 97892 35896 97894
rect 4220 97402 4276 97404
rect 4300 97402 4356 97404
rect 4380 97402 4436 97404
rect 4460 97402 4516 97404
rect 4220 97350 4266 97402
rect 4266 97350 4276 97402
rect 4300 97350 4330 97402
rect 4330 97350 4342 97402
rect 4342 97350 4356 97402
rect 4380 97350 4394 97402
rect 4394 97350 4406 97402
rect 4406 97350 4436 97402
rect 4460 97350 4470 97402
rect 4470 97350 4516 97402
rect 4220 97348 4276 97350
rect 4300 97348 4356 97350
rect 4380 97348 4436 97350
rect 4460 97348 4516 97350
rect 34940 97402 34996 97404
rect 35020 97402 35076 97404
rect 35100 97402 35156 97404
rect 35180 97402 35236 97404
rect 34940 97350 34986 97402
rect 34986 97350 34996 97402
rect 35020 97350 35050 97402
rect 35050 97350 35062 97402
rect 35062 97350 35076 97402
rect 35100 97350 35114 97402
rect 35114 97350 35126 97402
rect 35126 97350 35156 97402
rect 35180 97350 35190 97402
rect 35190 97350 35236 97402
rect 34940 97348 34996 97350
rect 35020 97348 35076 97350
rect 35100 97348 35156 97350
rect 35180 97348 35236 97350
rect 4880 96858 4936 96860
rect 4960 96858 5016 96860
rect 5040 96858 5096 96860
rect 5120 96858 5176 96860
rect 4880 96806 4926 96858
rect 4926 96806 4936 96858
rect 4960 96806 4990 96858
rect 4990 96806 5002 96858
rect 5002 96806 5016 96858
rect 5040 96806 5054 96858
rect 5054 96806 5066 96858
rect 5066 96806 5096 96858
rect 5120 96806 5130 96858
rect 5130 96806 5176 96858
rect 4880 96804 4936 96806
rect 4960 96804 5016 96806
rect 5040 96804 5096 96806
rect 5120 96804 5176 96806
rect 35600 96858 35656 96860
rect 35680 96858 35736 96860
rect 35760 96858 35816 96860
rect 35840 96858 35896 96860
rect 35600 96806 35646 96858
rect 35646 96806 35656 96858
rect 35680 96806 35710 96858
rect 35710 96806 35722 96858
rect 35722 96806 35736 96858
rect 35760 96806 35774 96858
rect 35774 96806 35786 96858
rect 35786 96806 35816 96858
rect 35840 96806 35850 96858
rect 35850 96806 35896 96858
rect 35600 96804 35656 96806
rect 35680 96804 35736 96806
rect 35760 96804 35816 96806
rect 35840 96804 35896 96806
rect 4220 96314 4276 96316
rect 4300 96314 4356 96316
rect 4380 96314 4436 96316
rect 4460 96314 4516 96316
rect 4220 96262 4266 96314
rect 4266 96262 4276 96314
rect 4300 96262 4330 96314
rect 4330 96262 4342 96314
rect 4342 96262 4356 96314
rect 4380 96262 4394 96314
rect 4394 96262 4406 96314
rect 4406 96262 4436 96314
rect 4460 96262 4470 96314
rect 4470 96262 4516 96314
rect 4220 96260 4276 96262
rect 4300 96260 4356 96262
rect 4380 96260 4436 96262
rect 4460 96260 4516 96262
rect 34940 96314 34996 96316
rect 35020 96314 35076 96316
rect 35100 96314 35156 96316
rect 35180 96314 35236 96316
rect 34940 96262 34986 96314
rect 34986 96262 34996 96314
rect 35020 96262 35050 96314
rect 35050 96262 35062 96314
rect 35062 96262 35076 96314
rect 35100 96262 35114 96314
rect 35114 96262 35126 96314
rect 35126 96262 35156 96314
rect 35180 96262 35190 96314
rect 35190 96262 35236 96314
rect 34940 96260 34996 96262
rect 35020 96260 35076 96262
rect 35100 96260 35156 96262
rect 35180 96260 35236 96262
rect 4880 95770 4936 95772
rect 4960 95770 5016 95772
rect 5040 95770 5096 95772
rect 5120 95770 5176 95772
rect 4880 95718 4926 95770
rect 4926 95718 4936 95770
rect 4960 95718 4990 95770
rect 4990 95718 5002 95770
rect 5002 95718 5016 95770
rect 5040 95718 5054 95770
rect 5054 95718 5066 95770
rect 5066 95718 5096 95770
rect 5120 95718 5130 95770
rect 5130 95718 5176 95770
rect 4880 95716 4936 95718
rect 4960 95716 5016 95718
rect 5040 95716 5096 95718
rect 5120 95716 5176 95718
rect 35600 95770 35656 95772
rect 35680 95770 35736 95772
rect 35760 95770 35816 95772
rect 35840 95770 35896 95772
rect 35600 95718 35646 95770
rect 35646 95718 35656 95770
rect 35680 95718 35710 95770
rect 35710 95718 35722 95770
rect 35722 95718 35736 95770
rect 35760 95718 35774 95770
rect 35774 95718 35786 95770
rect 35786 95718 35816 95770
rect 35840 95718 35850 95770
rect 35850 95718 35896 95770
rect 35600 95716 35656 95718
rect 35680 95716 35736 95718
rect 35760 95716 35816 95718
rect 35840 95716 35896 95718
rect 4220 95226 4276 95228
rect 4300 95226 4356 95228
rect 4380 95226 4436 95228
rect 4460 95226 4516 95228
rect 4220 95174 4266 95226
rect 4266 95174 4276 95226
rect 4300 95174 4330 95226
rect 4330 95174 4342 95226
rect 4342 95174 4356 95226
rect 4380 95174 4394 95226
rect 4394 95174 4406 95226
rect 4406 95174 4436 95226
rect 4460 95174 4470 95226
rect 4470 95174 4516 95226
rect 4220 95172 4276 95174
rect 4300 95172 4356 95174
rect 4380 95172 4436 95174
rect 4460 95172 4516 95174
rect 34940 95226 34996 95228
rect 35020 95226 35076 95228
rect 35100 95226 35156 95228
rect 35180 95226 35236 95228
rect 34940 95174 34986 95226
rect 34986 95174 34996 95226
rect 35020 95174 35050 95226
rect 35050 95174 35062 95226
rect 35062 95174 35076 95226
rect 35100 95174 35114 95226
rect 35114 95174 35126 95226
rect 35126 95174 35156 95226
rect 35180 95174 35190 95226
rect 35190 95174 35236 95226
rect 34940 95172 34996 95174
rect 35020 95172 35076 95174
rect 35100 95172 35156 95174
rect 35180 95172 35236 95174
rect 4880 94682 4936 94684
rect 4960 94682 5016 94684
rect 5040 94682 5096 94684
rect 5120 94682 5176 94684
rect 4880 94630 4926 94682
rect 4926 94630 4936 94682
rect 4960 94630 4990 94682
rect 4990 94630 5002 94682
rect 5002 94630 5016 94682
rect 5040 94630 5054 94682
rect 5054 94630 5066 94682
rect 5066 94630 5096 94682
rect 5120 94630 5130 94682
rect 5130 94630 5176 94682
rect 4880 94628 4936 94630
rect 4960 94628 5016 94630
rect 5040 94628 5096 94630
rect 5120 94628 5176 94630
rect 35600 94682 35656 94684
rect 35680 94682 35736 94684
rect 35760 94682 35816 94684
rect 35840 94682 35896 94684
rect 35600 94630 35646 94682
rect 35646 94630 35656 94682
rect 35680 94630 35710 94682
rect 35710 94630 35722 94682
rect 35722 94630 35736 94682
rect 35760 94630 35774 94682
rect 35774 94630 35786 94682
rect 35786 94630 35816 94682
rect 35840 94630 35850 94682
rect 35850 94630 35896 94682
rect 35600 94628 35656 94630
rect 35680 94628 35736 94630
rect 35760 94628 35816 94630
rect 35840 94628 35896 94630
rect 4220 94138 4276 94140
rect 4300 94138 4356 94140
rect 4380 94138 4436 94140
rect 4460 94138 4516 94140
rect 4220 94086 4266 94138
rect 4266 94086 4276 94138
rect 4300 94086 4330 94138
rect 4330 94086 4342 94138
rect 4342 94086 4356 94138
rect 4380 94086 4394 94138
rect 4394 94086 4406 94138
rect 4406 94086 4436 94138
rect 4460 94086 4470 94138
rect 4470 94086 4516 94138
rect 4220 94084 4276 94086
rect 4300 94084 4356 94086
rect 4380 94084 4436 94086
rect 4460 94084 4516 94086
rect 34940 94138 34996 94140
rect 35020 94138 35076 94140
rect 35100 94138 35156 94140
rect 35180 94138 35236 94140
rect 34940 94086 34986 94138
rect 34986 94086 34996 94138
rect 35020 94086 35050 94138
rect 35050 94086 35062 94138
rect 35062 94086 35076 94138
rect 35100 94086 35114 94138
rect 35114 94086 35126 94138
rect 35126 94086 35156 94138
rect 35180 94086 35190 94138
rect 35190 94086 35236 94138
rect 34940 94084 34996 94086
rect 35020 94084 35076 94086
rect 35100 94084 35156 94086
rect 35180 94084 35236 94086
rect 4880 93594 4936 93596
rect 4960 93594 5016 93596
rect 5040 93594 5096 93596
rect 5120 93594 5176 93596
rect 4880 93542 4926 93594
rect 4926 93542 4936 93594
rect 4960 93542 4990 93594
rect 4990 93542 5002 93594
rect 5002 93542 5016 93594
rect 5040 93542 5054 93594
rect 5054 93542 5066 93594
rect 5066 93542 5096 93594
rect 5120 93542 5130 93594
rect 5130 93542 5176 93594
rect 4880 93540 4936 93542
rect 4960 93540 5016 93542
rect 5040 93540 5096 93542
rect 5120 93540 5176 93542
rect 35600 93594 35656 93596
rect 35680 93594 35736 93596
rect 35760 93594 35816 93596
rect 35840 93594 35896 93596
rect 35600 93542 35646 93594
rect 35646 93542 35656 93594
rect 35680 93542 35710 93594
rect 35710 93542 35722 93594
rect 35722 93542 35736 93594
rect 35760 93542 35774 93594
rect 35774 93542 35786 93594
rect 35786 93542 35816 93594
rect 35840 93542 35850 93594
rect 35850 93542 35896 93594
rect 35600 93540 35656 93542
rect 35680 93540 35736 93542
rect 35760 93540 35816 93542
rect 35840 93540 35896 93542
rect 4220 93050 4276 93052
rect 4300 93050 4356 93052
rect 4380 93050 4436 93052
rect 4460 93050 4516 93052
rect 4220 92998 4266 93050
rect 4266 92998 4276 93050
rect 4300 92998 4330 93050
rect 4330 92998 4342 93050
rect 4342 92998 4356 93050
rect 4380 92998 4394 93050
rect 4394 92998 4406 93050
rect 4406 92998 4436 93050
rect 4460 92998 4470 93050
rect 4470 92998 4516 93050
rect 4220 92996 4276 92998
rect 4300 92996 4356 92998
rect 4380 92996 4436 92998
rect 4460 92996 4516 92998
rect 34940 93050 34996 93052
rect 35020 93050 35076 93052
rect 35100 93050 35156 93052
rect 35180 93050 35236 93052
rect 34940 92998 34986 93050
rect 34986 92998 34996 93050
rect 35020 92998 35050 93050
rect 35050 92998 35062 93050
rect 35062 92998 35076 93050
rect 35100 92998 35114 93050
rect 35114 92998 35126 93050
rect 35126 92998 35156 93050
rect 35180 92998 35190 93050
rect 35190 92998 35236 93050
rect 34940 92996 34996 92998
rect 35020 92996 35076 92998
rect 35100 92996 35156 92998
rect 35180 92996 35236 92998
rect 4880 92506 4936 92508
rect 4960 92506 5016 92508
rect 5040 92506 5096 92508
rect 5120 92506 5176 92508
rect 4880 92454 4926 92506
rect 4926 92454 4936 92506
rect 4960 92454 4990 92506
rect 4990 92454 5002 92506
rect 5002 92454 5016 92506
rect 5040 92454 5054 92506
rect 5054 92454 5066 92506
rect 5066 92454 5096 92506
rect 5120 92454 5130 92506
rect 5130 92454 5176 92506
rect 4880 92452 4936 92454
rect 4960 92452 5016 92454
rect 5040 92452 5096 92454
rect 5120 92452 5176 92454
rect 35600 92506 35656 92508
rect 35680 92506 35736 92508
rect 35760 92506 35816 92508
rect 35840 92506 35896 92508
rect 35600 92454 35646 92506
rect 35646 92454 35656 92506
rect 35680 92454 35710 92506
rect 35710 92454 35722 92506
rect 35722 92454 35736 92506
rect 35760 92454 35774 92506
rect 35774 92454 35786 92506
rect 35786 92454 35816 92506
rect 35840 92454 35850 92506
rect 35850 92454 35896 92506
rect 35600 92452 35656 92454
rect 35680 92452 35736 92454
rect 35760 92452 35816 92454
rect 35840 92452 35896 92454
rect 4220 91962 4276 91964
rect 4300 91962 4356 91964
rect 4380 91962 4436 91964
rect 4460 91962 4516 91964
rect 4220 91910 4266 91962
rect 4266 91910 4276 91962
rect 4300 91910 4330 91962
rect 4330 91910 4342 91962
rect 4342 91910 4356 91962
rect 4380 91910 4394 91962
rect 4394 91910 4406 91962
rect 4406 91910 4436 91962
rect 4460 91910 4470 91962
rect 4470 91910 4516 91962
rect 4220 91908 4276 91910
rect 4300 91908 4356 91910
rect 4380 91908 4436 91910
rect 4460 91908 4516 91910
rect 34940 91962 34996 91964
rect 35020 91962 35076 91964
rect 35100 91962 35156 91964
rect 35180 91962 35236 91964
rect 34940 91910 34986 91962
rect 34986 91910 34996 91962
rect 35020 91910 35050 91962
rect 35050 91910 35062 91962
rect 35062 91910 35076 91962
rect 35100 91910 35114 91962
rect 35114 91910 35126 91962
rect 35126 91910 35156 91962
rect 35180 91910 35190 91962
rect 35190 91910 35236 91962
rect 34940 91908 34996 91910
rect 35020 91908 35076 91910
rect 35100 91908 35156 91910
rect 35180 91908 35236 91910
rect 4880 91418 4936 91420
rect 4960 91418 5016 91420
rect 5040 91418 5096 91420
rect 5120 91418 5176 91420
rect 4880 91366 4926 91418
rect 4926 91366 4936 91418
rect 4960 91366 4990 91418
rect 4990 91366 5002 91418
rect 5002 91366 5016 91418
rect 5040 91366 5054 91418
rect 5054 91366 5066 91418
rect 5066 91366 5096 91418
rect 5120 91366 5130 91418
rect 5130 91366 5176 91418
rect 4880 91364 4936 91366
rect 4960 91364 5016 91366
rect 5040 91364 5096 91366
rect 5120 91364 5176 91366
rect 35600 91418 35656 91420
rect 35680 91418 35736 91420
rect 35760 91418 35816 91420
rect 35840 91418 35896 91420
rect 35600 91366 35646 91418
rect 35646 91366 35656 91418
rect 35680 91366 35710 91418
rect 35710 91366 35722 91418
rect 35722 91366 35736 91418
rect 35760 91366 35774 91418
rect 35774 91366 35786 91418
rect 35786 91366 35816 91418
rect 35840 91366 35850 91418
rect 35850 91366 35896 91418
rect 35600 91364 35656 91366
rect 35680 91364 35736 91366
rect 35760 91364 35816 91366
rect 35840 91364 35896 91366
rect 4220 90874 4276 90876
rect 4300 90874 4356 90876
rect 4380 90874 4436 90876
rect 4460 90874 4516 90876
rect 4220 90822 4266 90874
rect 4266 90822 4276 90874
rect 4300 90822 4330 90874
rect 4330 90822 4342 90874
rect 4342 90822 4356 90874
rect 4380 90822 4394 90874
rect 4394 90822 4406 90874
rect 4406 90822 4436 90874
rect 4460 90822 4470 90874
rect 4470 90822 4516 90874
rect 4220 90820 4276 90822
rect 4300 90820 4356 90822
rect 4380 90820 4436 90822
rect 4460 90820 4516 90822
rect 34940 90874 34996 90876
rect 35020 90874 35076 90876
rect 35100 90874 35156 90876
rect 35180 90874 35236 90876
rect 34940 90822 34986 90874
rect 34986 90822 34996 90874
rect 35020 90822 35050 90874
rect 35050 90822 35062 90874
rect 35062 90822 35076 90874
rect 35100 90822 35114 90874
rect 35114 90822 35126 90874
rect 35126 90822 35156 90874
rect 35180 90822 35190 90874
rect 35190 90822 35236 90874
rect 34940 90820 34996 90822
rect 35020 90820 35076 90822
rect 35100 90820 35156 90822
rect 35180 90820 35236 90822
rect 4880 90330 4936 90332
rect 4960 90330 5016 90332
rect 5040 90330 5096 90332
rect 5120 90330 5176 90332
rect 4880 90278 4926 90330
rect 4926 90278 4936 90330
rect 4960 90278 4990 90330
rect 4990 90278 5002 90330
rect 5002 90278 5016 90330
rect 5040 90278 5054 90330
rect 5054 90278 5066 90330
rect 5066 90278 5096 90330
rect 5120 90278 5130 90330
rect 5130 90278 5176 90330
rect 4880 90276 4936 90278
rect 4960 90276 5016 90278
rect 5040 90276 5096 90278
rect 5120 90276 5176 90278
rect 35600 90330 35656 90332
rect 35680 90330 35736 90332
rect 35760 90330 35816 90332
rect 35840 90330 35896 90332
rect 35600 90278 35646 90330
rect 35646 90278 35656 90330
rect 35680 90278 35710 90330
rect 35710 90278 35722 90330
rect 35722 90278 35736 90330
rect 35760 90278 35774 90330
rect 35774 90278 35786 90330
rect 35786 90278 35816 90330
rect 35840 90278 35850 90330
rect 35850 90278 35896 90330
rect 35600 90276 35656 90278
rect 35680 90276 35736 90278
rect 35760 90276 35816 90278
rect 35840 90276 35896 90278
rect 4220 89786 4276 89788
rect 4300 89786 4356 89788
rect 4380 89786 4436 89788
rect 4460 89786 4516 89788
rect 4220 89734 4266 89786
rect 4266 89734 4276 89786
rect 4300 89734 4330 89786
rect 4330 89734 4342 89786
rect 4342 89734 4356 89786
rect 4380 89734 4394 89786
rect 4394 89734 4406 89786
rect 4406 89734 4436 89786
rect 4460 89734 4470 89786
rect 4470 89734 4516 89786
rect 4220 89732 4276 89734
rect 4300 89732 4356 89734
rect 4380 89732 4436 89734
rect 4460 89732 4516 89734
rect 34940 89786 34996 89788
rect 35020 89786 35076 89788
rect 35100 89786 35156 89788
rect 35180 89786 35236 89788
rect 34940 89734 34986 89786
rect 34986 89734 34996 89786
rect 35020 89734 35050 89786
rect 35050 89734 35062 89786
rect 35062 89734 35076 89786
rect 35100 89734 35114 89786
rect 35114 89734 35126 89786
rect 35126 89734 35156 89786
rect 35180 89734 35190 89786
rect 35190 89734 35236 89786
rect 34940 89732 34996 89734
rect 35020 89732 35076 89734
rect 35100 89732 35156 89734
rect 35180 89732 35236 89734
rect 4880 89242 4936 89244
rect 4960 89242 5016 89244
rect 5040 89242 5096 89244
rect 5120 89242 5176 89244
rect 4880 89190 4926 89242
rect 4926 89190 4936 89242
rect 4960 89190 4990 89242
rect 4990 89190 5002 89242
rect 5002 89190 5016 89242
rect 5040 89190 5054 89242
rect 5054 89190 5066 89242
rect 5066 89190 5096 89242
rect 5120 89190 5130 89242
rect 5130 89190 5176 89242
rect 4880 89188 4936 89190
rect 4960 89188 5016 89190
rect 5040 89188 5096 89190
rect 5120 89188 5176 89190
rect 35600 89242 35656 89244
rect 35680 89242 35736 89244
rect 35760 89242 35816 89244
rect 35840 89242 35896 89244
rect 35600 89190 35646 89242
rect 35646 89190 35656 89242
rect 35680 89190 35710 89242
rect 35710 89190 35722 89242
rect 35722 89190 35736 89242
rect 35760 89190 35774 89242
rect 35774 89190 35786 89242
rect 35786 89190 35816 89242
rect 35840 89190 35850 89242
rect 35850 89190 35896 89242
rect 35600 89188 35656 89190
rect 35680 89188 35736 89190
rect 35760 89188 35816 89190
rect 35840 89188 35896 89190
rect 4220 88698 4276 88700
rect 4300 88698 4356 88700
rect 4380 88698 4436 88700
rect 4460 88698 4516 88700
rect 4220 88646 4266 88698
rect 4266 88646 4276 88698
rect 4300 88646 4330 88698
rect 4330 88646 4342 88698
rect 4342 88646 4356 88698
rect 4380 88646 4394 88698
rect 4394 88646 4406 88698
rect 4406 88646 4436 88698
rect 4460 88646 4470 88698
rect 4470 88646 4516 88698
rect 4220 88644 4276 88646
rect 4300 88644 4356 88646
rect 4380 88644 4436 88646
rect 4460 88644 4516 88646
rect 34940 88698 34996 88700
rect 35020 88698 35076 88700
rect 35100 88698 35156 88700
rect 35180 88698 35236 88700
rect 34940 88646 34986 88698
rect 34986 88646 34996 88698
rect 35020 88646 35050 88698
rect 35050 88646 35062 88698
rect 35062 88646 35076 88698
rect 35100 88646 35114 88698
rect 35114 88646 35126 88698
rect 35126 88646 35156 88698
rect 35180 88646 35190 88698
rect 35190 88646 35236 88698
rect 34940 88644 34996 88646
rect 35020 88644 35076 88646
rect 35100 88644 35156 88646
rect 35180 88644 35236 88646
rect 4880 88154 4936 88156
rect 4960 88154 5016 88156
rect 5040 88154 5096 88156
rect 5120 88154 5176 88156
rect 4880 88102 4926 88154
rect 4926 88102 4936 88154
rect 4960 88102 4990 88154
rect 4990 88102 5002 88154
rect 5002 88102 5016 88154
rect 5040 88102 5054 88154
rect 5054 88102 5066 88154
rect 5066 88102 5096 88154
rect 5120 88102 5130 88154
rect 5130 88102 5176 88154
rect 4880 88100 4936 88102
rect 4960 88100 5016 88102
rect 5040 88100 5096 88102
rect 5120 88100 5176 88102
rect 35600 88154 35656 88156
rect 35680 88154 35736 88156
rect 35760 88154 35816 88156
rect 35840 88154 35896 88156
rect 35600 88102 35646 88154
rect 35646 88102 35656 88154
rect 35680 88102 35710 88154
rect 35710 88102 35722 88154
rect 35722 88102 35736 88154
rect 35760 88102 35774 88154
rect 35774 88102 35786 88154
rect 35786 88102 35816 88154
rect 35840 88102 35850 88154
rect 35850 88102 35896 88154
rect 35600 88100 35656 88102
rect 35680 88100 35736 88102
rect 35760 88100 35816 88102
rect 35840 88100 35896 88102
rect 4220 87610 4276 87612
rect 4300 87610 4356 87612
rect 4380 87610 4436 87612
rect 4460 87610 4516 87612
rect 4220 87558 4266 87610
rect 4266 87558 4276 87610
rect 4300 87558 4330 87610
rect 4330 87558 4342 87610
rect 4342 87558 4356 87610
rect 4380 87558 4394 87610
rect 4394 87558 4406 87610
rect 4406 87558 4436 87610
rect 4460 87558 4470 87610
rect 4470 87558 4516 87610
rect 4220 87556 4276 87558
rect 4300 87556 4356 87558
rect 4380 87556 4436 87558
rect 4460 87556 4516 87558
rect 34940 87610 34996 87612
rect 35020 87610 35076 87612
rect 35100 87610 35156 87612
rect 35180 87610 35236 87612
rect 34940 87558 34986 87610
rect 34986 87558 34996 87610
rect 35020 87558 35050 87610
rect 35050 87558 35062 87610
rect 35062 87558 35076 87610
rect 35100 87558 35114 87610
rect 35114 87558 35126 87610
rect 35126 87558 35156 87610
rect 35180 87558 35190 87610
rect 35190 87558 35236 87610
rect 34940 87556 34996 87558
rect 35020 87556 35076 87558
rect 35100 87556 35156 87558
rect 35180 87556 35236 87558
rect 4880 87066 4936 87068
rect 4960 87066 5016 87068
rect 5040 87066 5096 87068
rect 5120 87066 5176 87068
rect 4880 87014 4926 87066
rect 4926 87014 4936 87066
rect 4960 87014 4990 87066
rect 4990 87014 5002 87066
rect 5002 87014 5016 87066
rect 5040 87014 5054 87066
rect 5054 87014 5066 87066
rect 5066 87014 5096 87066
rect 5120 87014 5130 87066
rect 5130 87014 5176 87066
rect 4880 87012 4936 87014
rect 4960 87012 5016 87014
rect 5040 87012 5096 87014
rect 5120 87012 5176 87014
rect 35600 87066 35656 87068
rect 35680 87066 35736 87068
rect 35760 87066 35816 87068
rect 35840 87066 35896 87068
rect 35600 87014 35646 87066
rect 35646 87014 35656 87066
rect 35680 87014 35710 87066
rect 35710 87014 35722 87066
rect 35722 87014 35736 87066
rect 35760 87014 35774 87066
rect 35774 87014 35786 87066
rect 35786 87014 35816 87066
rect 35840 87014 35850 87066
rect 35850 87014 35896 87066
rect 35600 87012 35656 87014
rect 35680 87012 35736 87014
rect 35760 87012 35816 87014
rect 35840 87012 35896 87014
rect 4220 86522 4276 86524
rect 4300 86522 4356 86524
rect 4380 86522 4436 86524
rect 4460 86522 4516 86524
rect 4220 86470 4266 86522
rect 4266 86470 4276 86522
rect 4300 86470 4330 86522
rect 4330 86470 4342 86522
rect 4342 86470 4356 86522
rect 4380 86470 4394 86522
rect 4394 86470 4406 86522
rect 4406 86470 4436 86522
rect 4460 86470 4470 86522
rect 4470 86470 4516 86522
rect 4220 86468 4276 86470
rect 4300 86468 4356 86470
rect 4380 86468 4436 86470
rect 4460 86468 4516 86470
rect 34940 86522 34996 86524
rect 35020 86522 35076 86524
rect 35100 86522 35156 86524
rect 35180 86522 35236 86524
rect 34940 86470 34986 86522
rect 34986 86470 34996 86522
rect 35020 86470 35050 86522
rect 35050 86470 35062 86522
rect 35062 86470 35076 86522
rect 35100 86470 35114 86522
rect 35114 86470 35126 86522
rect 35126 86470 35156 86522
rect 35180 86470 35190 86522
rect 35190 86470 35236 86522
rect 34940 86468 34996 86470
rect 35020 86468 35076 86470
rect 35100 86468 35156 86470
rect 35180 86468 35236 86470
rect 4880 85978 4936 85980
rect 4960 85978 5016 85980
rect 5040 85978 5096 85980
rect 5120 85978 5176 85980
rect 4880 85926 4926 85978
rect 4926 85926 4936 85978
rect 4960 85926 4990 85978
rect 4990 85926 5002 85978
rect 5002 85926 5016 85978
rect 5040 85926 5054 85978
rect 5054 85926 5066 85978
rect 5066 85926 5096 85978
rect 5120 85926 5130 85978
rect 5130 85926 5176 85978
rect 4880 85924 4936 85926
rect 4960 85924 5016 85926
rect 5040 85924 5096 85926
rect 5120 85924 5176 85926
rect 35600 85978 35656 85980
rect 35680 85978 35736 85980
rect 35760 85978 35816 85980
rect 35840 85978 35896 85980
rect 35600 85926 35646 85978
rect 35646 85926 35656 85978
rect 35680 85926 35710 85978
rect 35710 85926 35722 85978
rect 35722 85926 35736 85978
rect 35760 85926 35774 85978
rect 35774 85926 35786 85978
rect 35786 85926 35816 85978
rect 35840 85926 35850 85978
rect 35850 85926 35896 85978
rect 35600 85924 35656 85926
rect 35680 85924 35736 85926
rect 35760 85924 35816 85926
rect 35840 85924 35896 85926
rect 4220 85434 4276 85436
rect 4300 85434 4356 85436
rect 4380 85434 4436 85436
rect 4460 85434 4516 85436
rect 4220 85382 4266 85434
rect 4266 85382 4276 85434
rect 4300 85382 4330 85434
rect 4330 85382 4342 85434
rect 4342 85382 4356 85434
rect 4380 85382 4394 85434
rect 4394 85382 4406 85434
rect 4406 85382 4436 85434
rect 4460 85382 4470 85434
rect 4470 85382 4516 85434
rect 4220 85380 4276 85382
rect 4300 85380 4356 85382
rect 4380 85380 4436 85382
rect 4460 85380 4516 85382
rect 34940 85434 34996 85436
rect 35020 85434 35076 85436
rect 35100 85434 35156 85436
rect 35180 85434 35236 85436
rect 34940 85382 34986 85434
rect 34986 85382 34996 85434
rect 35020 85382 35050 85434
rect 35050 85382 35062 85434
rect 35062 85382 35076 85434
rect 35100 85382 35114 85434
rect 35114 85382 35126 85434
rect 35126 85382 35156 85434
rect 35180 85382 35190 85434
rect 35190 85382 35236 85434
rect 34940 85380 34996 85382
rect 35020 85380 35076 85382
rect 35100 85380 35156 85382
rect 35180 85380 35236 85382
rect 4880 84890 4936 84892
rect 4960 84890 5016 84892
rect 5040 84890 5096 84892
rect 5120 84890 5176 84892
rect 4880 84838 4926 84890
rect 4926 84838 4936 84890
rect 4960 84838 4990 84890
rect 4990 84838 5002 84890
rect 5002 84838 5016 84890
rect 5040 84838 5054 84890
rect 5054 84838 5066 84890
rect 5066 84838 5096 84890
rect 5120 84838 5130 84890
rect 5130 84838 5176 84890
rect 4880 84836 4936 84838
rect 4960 84836 5016 84838
rect 5040 84836 5096 84838
rect 5120 84836 5176 84838
rect 35600 84890 35656 84892
rect 35680 84890 35736 84892
rect 35760 84890 35816 84892
rect 35840 84890 35896 84892
rect 35600 84838 35646 84890
rect 35646 84838 35656 84890
rect 35680 84838 35710 84890
rect 35710 84838 35722 84890
rect 35722 84838 35736 84890
rect 35760 84838 35774 84890
rect 35774 84838 35786 84890
rect 35786 84838 35816 84890
rect 35840 84838 35850 84890
rect 35850 84838 35896 84890
rect 35600 84836 35656 84838
rect 35680 84836 35736 84838
rect 35760 84836 35816 84838
rect 35840 84836 35896 84838
rect 4220 84346 4276 84348
rect 4300 84346 4356 84348
rect 4380 84346 4436 84348
rect 4460 84346 4516 84348
rect 4220 84294 4266 84346
rect 4266 84294 4276 84346
rect 4300 84294 4330 84346
rect 4330 84294 4342 84346
rect 4342 84294 4356 84346
rect 4380 84294 4394 84346
rect 4394 84294 4406 84346
rect 4406 84294 4436 84346
rect 4460 84294 4470 84346
rect 4470 84294 4516 84346
rect 4220 84292 4276 84294
rect 4300 84292 4356 84294
rect 4380 84292 4436 84294
rect 4460 84292 4516 84294
rect 34940 84346 34996 84348
rect 35020 84346 35076 84348
rect 35100 84346 35156 84348
rect 35180 84346 35236 84348
rect 34940 84294 34986 84346
rect 34986 84294 34996 84346
rect 35020 84294 35050 84346
rect 35050 84294 35062 84346
rect 35062 84294 35076 84346
rect 35100 84294 35114 84346
rect 35114 84294 35126 84346
rect 35126 84294 35156 84346
rect 35180 84294 35190 84346
rect 35190 84294 35236 84346
rect 34940 84292 34996 84294
rect 35020 84292 35076 84294
rect 35100 84292 35156 84294
rect 35180 84292 35236 84294
rect 4880 83802 4936 83804
rect 4960 83802 5016 83804
rect 5040 83802 5096 83804
rect 5120 83802 5176 83804
rect 4880 83750 4926 83802
rect 4926 83750 4936 83802
rect 4960 83750 4990 83802
rect 4990 83750 5002 83802
rect 5002 83750 5016 83802
rect 5040 83750 5054 83802
rect 5054 83750 5066 83802
rect 5066 83750 5096 83802
rect 5120 83750 5130 83802
rect 5130 83750 5176 83802
rect 4880 83748 4936 83750
rect 4960 83748 5016 83750
rect 5040 83748 5096 83750
rect 5120 83748 5176 83750
rect 35600 83802 35656 83804
rect 35680 83802 35736 83804
rect 35760 83802 35816 83804
rect 35840 83802 35896 83804
rect 35600 83750 35646 83802
rect 35646 83750 35656 83802
rect 35680 83750 35710 83802
rect 35710 83750 35722 83802
rect 35722 83750 35736 83802
rect 35760 83750 35774 83802
rect 35774 83750 35786 83802
rect 35786 83750 35816 83802
rect 35840 83750 35850 83802
rect 35850 83750 35896 83802
rect 35600 83748 35656 83750
rect 35680 83748 35736 83750
rect 35760 83748 35816 83750
rect 35840 83748 35896 83750
rect 4220 83258 4276 83260
rect 4300 83258 4356 83260
rect 4380 83258 4436 83260
rect 4460 83258 4516 83260
rect 4220 83206 4266 83258
rect 4266 83206 4276 83258
rect 4300 83206 4330 83258
rect 4330 83206 4342 83258
rect 4342 83206 4356 83258
rect 4380 83206 4394 83258
rect 4394 83206 4406 83258
rect 4406 83206 4436 83258
rect 4460 83206 4470 83258
rect 4470 83206 4516 83258
rect 4220 83204 4276 83206
rect 4300 83204 4356 83206
rect 4380 83204 4436 83206
rect 4460 83204 4516 83206
rect 34940 83258 34996 83260
rect 35020 83258 35076 83260
rect 35100 83258 35156 83260
rect 35180 83258 35236 83260
rect 34940 83206 34986 83258
rect 34986 83206 34996 83258
rect 35020 83206 35050 83258
rect 35050 83206 35062 83258
rect 35062 83206 35076 83258
rect 35100 83206 35114 83258
rect 35114 83206 35126 83258
rect 35126 83206 35156 83258
rect 35180 83206 35190 83258
rect 35190 83206 35236 83258
rect 34940 83204 34996 83206
rect 35020 83204 35076 83206
rect 35100 83204 35156 83206
rect 35180 83204 35236 83206
rect 4880 82714 4936 82716
rect 4960 82714 5016 82716
rect 5040 82714 5096 82716
rect 5120 82714 5176 82716
rect 4880 82662 4926 82714
rect 4926 82662 4936 82714
rect 4960 82662 4990 82714
rect 4990 82662 5002 82714
rect 5002 82662 5016 82714
rect 5040 82662 5054 82714
rect 5054 82662 5066 82714
rect 5066 82662 5096 82714
rect 5120 82662 5130 82714
rect 5130 82662 5176 82714
rect 4880 82660 4936 82662
rect 4960 82660 5016 82662
rect 5040 82660 5096 82662
rect 5120 82660 5176 82662
rect 35600 82714 35656 82716
rect 35680 82714 35736 82716
rect 35760 82714 35816 82716
rect 35840 82714 35896 82716
rect 35600 82662 35646 82714
rect 35646 82662 35656 82714
rect 35680 82662 35710 82714
rect 35710 82662 35722 82714
rect 35722 82662 35736 82714
rect 35760 82662 35774 82714
rect 35774 82662 35786 82714
rect 35786 82662 35816 82714
rect 35840 82662 35850 82714
rect 35850 82662 35896 82714
rect 35600 82660 35656 82662
rect 35680 82660 35736 82662
rect 35760 82660 35816 82662
rect 35840 82660 35896 82662
rect 4220 82170 4276 82172
rect 4300 82170 4356 82172
rect 4380 82170 4436 82172
rect 4460 82170 4516 82172
rect 4220 82118 4266 82170
rect 4266 82118 4276 82170
rect 4300 82118 4330 82170
rect 4330 82118 4342 82170
rect 4342 82118 4356 82170
rect 4380 82118 4394 82170
rect 4394 82118 4406 82170
rect 4406 82118 4436 82170
rect 4460 82118 4470 82170
rect 4470 82118 4516 82170
rect 4220 82116 4276 82118
rect 4300 82116 4356 82118
rect 4380 82116 4436 82118
rect 4460 82116 4516 82118
rect 34940 82170 34996 82172
rect 35020 82170 35076 82172
rect 35100 82170 35156 82172
rect 35180 82170 35236 82172
rect 34940 82118 34986 82170
rect 34986 82118 34996 82170
rect 35020 82118 35050 82170
rect 35050 82118 35062 82170
rect 35062 82118 35076 82170
rect 35100 82118 35114 82170
rect 35114 82118 35126 82170
rect 35126 82118 35156 82170
rect 35180 82118 35190 82170
rect 35190 82118 35236 82170
rect 34940 82116 34996 82118
rect 35020 82116 35076 82118
rect 35100 82116 35156 82118
rect 35180 82116 35236 82118
rect 4880 81626 4936 81628
rect 4960 81626 5016 81628
rect 5040 81626 5096 81628
rect 5120 81626 5176 81628
rect 4880 81574 4926 81626
rect 4926 81574 4936 81626
rect 4960 81574 4990 81626
rect 4990 81574 5002 81626
rect 5002 81574 5016 81626
rect 5040 81574 5054 81626
rect 5054 81574 5066 81626
rect 5066 81574 5096 81626
rect 5120 81574 5130 81626
rect 5130 81574 5176 81626
rect 4880 81572 4936 81574
rect 4960 81572 5016 81574
rect 5040 81572 5096 81574
rect 5120 81572 5176 81574
rect 35600 81626 35656 81628
rect 35680 81626 35736 81628
rect 35760 81626 35816 81628
rect 35840 81626 35896 81628
rect 35600 81574 35646 81626
rect 35646 81574 35656 81626
rect 35680 81574 35710 81626
rect 35710 81574 35722 81626
rect 35722 81574 35736 81626
rect 35760 81574 35774 81626
rect 35774 81574 35786 81626
rect 35786 81574 35816 81626
rect 35840 81574 35850 81626
rect 35850 81574 35896 81626
rect 35600 81572 35656 81574
rect 35680 81572 35736 81574
rect 35760 81572 35816 81574
rect 35840 81572 35896 81574
rect 4220 81082 4276 81084
rect 4300 81082 4356 81084
rect 4380 81082 4436 81084
rect 4460 81082 4516 81084
rect 4220 81030 4266 81082
rect 4266 81030 4276 81082
rect 4300 81030 4330 81082
rect 4330 81030 4342 81082
rect 4342 81030 4356 81082
rect 4380 81030 4394 81082
rect 4394 81030 4406 81082
rect 4406 81030 4436 81082
rect 4460 81030 4470 81082
rect 4470 81030 4516 81082
rect 4220 81028 4276 81030
rect 4300 81028 4356 81030
rect 4380 81028 4436 81030
rect 4460 81028 4516 81030
rect 34940 81082 34996 81084
rect 35020 81082 35076 81084
rect 35100 81082 35156 81084
rect 35180 81082 35236 81084
rect 34940 81030 34986 81082
rect 34986 81030 34996 81082
rect 35020 81030 35050 81082
rect 35050 81030 35062 81082
rect 35062 81030 35076 81082
rect 35100 81030 35114 81082
rect 35114 81030 35126 81082
rect 35126 81030 35156 81082
rect 35180 81030 35190 81082
rect 35190 81030 35236 81082
rect 34940 81028 34996 81030
rect 35020 81028 35076 81030
rect 35100 81028 35156 81030
rect 35180 81028 35236 81030
rect 4880 80538 4936 80540
rect 4960 80538 5016 80540
rect 5040 80538 5096 80540
rect 5120 80538 5176 80540
rect 4880 80486 4926 80538
rect 4926 80486 4936 80538
rect 4960 80486 4990 80538
rect 4990 80486 5002 80538
rect 5002 80486 5016 80538
rect 5040 80486 5054 80538
rect 5054 80486 5066 80538
rect 5066 80486 5096 80538
rect 5120 80486 5130 80538
rect 5130 80486 5176 80538
rect 4880 80484 4936 80486
rect 4960 80484 5016 80486
rect 5040 80484 5096 80486
rect 5120 80484 5176 80486
rect 35600 80538 35656 80540
rect 35680 80538 35736 80540
rect 35760 80538 35816 80540
rect 35840 80538 35896 80540
rect 35600 80486 35646 80538
rect 35646 80486 35656 80538
rect 35680 80486 35710 80538
rect 35710 80486 35722 80538
rect 35722 80486 35736 80538
rect 35760 80486 35774 80538
rect 35774 80486 35786 80538
rect 35786 80486 35816 80538
rect 35840 80486 35850 80538
rect 35850 80486 35896 80538
rect 35600 80484 35656 80486
rect 35680 80484 35736 80486
rect 35760 80484 35816 80486
rect 35840 80484 35896 80486
rect 4220 79994 4276 79996
rect 4300 79994 4356 79996
rect 4380 79994 4436 79996
rect 4460 79994 4516 79996
rect 4220 79942 4266 79994
rect 4266 79942 4276 79994
rect 4300 79942 4330 79994
rect 4330 79942 4342 79994
rect 4342 79942 4356 79994
rect 4380 79942 4394 79994
rect 4394 79942 4406 79994
rect 4406 79942 4436 79994
rect 4460 79942 4470 79994
rect 4470 79942 4516 79994
rect 4220 79940 4276 79942
rect 4300 79940 4356 79942
rect 4380 79940 4436 79942
rect 4460 79940 4516 79942
rect 34940 79994 34996 79996
rect 35020 79994 35076 79996
rect 35100 79994 35156 79996
rect 35180 79994 35236 79996
rect 34940 79942 34986 79994
rect 34986 79942 34996 79994
rect 35020 79942 35050 79994
rect 35050 79942 35062 79994
rect 35062 79942 35076 79994
rect 35100 79942 35114 79994
rect 35114 79942 35126 79994
rect 35126 79942 35156 79994
rect 35180 79942 35190 79994
rect 35190 79942 35236 79994
rect 34940 79940 34996 79942
rect 35020 79940 35076 79942
rect 35100 79940 35156 79942
rect 35180 79940 35236 79942
rect 4880 79450 4936 79452
rect 4960 79450 5016 79452
rect 5040 79450 5096 79452
rect 5120 79450 5176 79452
rect 4880 79398 4926 79450
rect 4926 79398 4936 79450
rect 4960 79398 4990 79450
rect 4990 79398 5002 79450
rect 5002 79398 5016 79450
rect 5040 79398 5054 79450
rect 5054 79398 5066 79450
rect 5066 79398 5096 79450
rect 5120 79398 5130 79450
rect 5130 79398 5176 79450
rect 4880 79396 4936 79398
rect 4960 79396 5016 79398
rect 5040 79396 5096 79398
rect 5120 79396 5176 79398
rect 35600 79450 35656 79452
rect 35680 79450 35736 79452
rect 35760 79450 35816 79452
rect 35840 79450 35896 79452
rect 35600 79398 35646 79450
rect 35646 79398 35656 79450
rect 35680 79398 35710 79450
rect 35710 79398 35722 79450
rect 35722 79398 35736 79450
rect 35760 79398 35774 79450
rect 35774 79398 35786 79450
rect 35786 79398 35816 79450
rect 35840 79398 35850 79450
rect 35850 79398 35896 79450
rect 35600 79396 35656 79398
rect 35680 79396 35736 79398
rect 35760 79396 35816 79398
rect 35840 79396 35896 79398
rect 4220 78906 4276 78908
rect 4300 78906 4356 78908
rect 4380 78906 4436 78908
rect 4460 78906 4516 78908
rect 4220 78854 4266 78906
rect 4266 78854 4276 78906
rect 4300 78854 4330 78906
rect 4330 78854 4342 78906
rect 4342 78854 4356 78906
rect 4380 78854 4394 78906
rect 4394 78854 4406 78906
rect 4406 78854 4436 78906
rect 4460 78854 4470 78906
rect 4470 78854 4516 78906
rect 4220 78852 4276 78854
rect 4300 78852 4356 78854
rect 4380 78852 4436 78854
rect 4460 78852 4516 78854
rect 34940 78906 34996 78908
rect 35020 78906 35076 78908
rect 35100 78906 35156 78908
rect 35180 78906 35236 78908
rect 34940 78854 34986 78906
rect 34986 78854 34996 78906
rect 35020 78854 35050 78906
rect 35050 78854 35062 78906
rect 35062 78854 35076 78906
rect 35100 78854 35114 78906
rect 35114 78854 35126 78906
rect 35126 78854 35156 78906
rect 35180 78854 35190 78906
rect 35190 78854 35236 78906
rect 34940 78852 34996 78854
rect 35020 78852 35076 78854
rect 35100 78852 35156 78854
rect 35180 78852 35236 78854
rect 4880 78362 4936 78364
rect 4960 78362 5016 78364
rect 5040 78362 5096 78364
rect 5120 78362 5176 78364
rect 4880 78310 4926 78362
rect 4926 78310 4936 78362
rect 4960 78310 4990 78362
rect 4990 78310 5002 78362
rect 5002 78310 5016 78362
rect 5040 78310 5054 78362
rect 5054 78310 5066 78362
rect 5066 78310 5096 78362
rect 5120 78310 5130 78362
rect 5130 78310 5176 78362
rect 4880 78308 4936 78310
rect 4960 78308 5016 78310
rect 5040 78308 5096 78310
rect 5120 78308 5176 78310
rect 35600 78362 35656 78364
rect 35680 78362 35736 78364
rect 35760 78362 35816 78364
rect 35840 78362 35896 78364
rect 35600 78310 35646 78362
rect 35646 78310 35656 78362
rect 35680 78310 35710 78362
rect 35710 78310 35722 78362
rect 35722 78310 35736 78362
rect 35760 78310 35774 78362
rect 35774 78310 35786 78362
rect 35786 78310 35816 78362
rect 35840 78310 35850 78362
rect 35850 78310 35896 78362
rect 35600 78308 35656 78310
rect 35680 78308 35736 78310
rect 35760 78308 35816 78310
rect 35840 78308 35896 78310
rect 4220 77818 4276 77820
rect 4300 77818 4356 77820
rect 4380 77818 4436 77820
rect 4460 77818 4516 77820
rect 4220 77766 4266 77818
rect 4266 77766 4276 77818
rect 4300 77766 4330 77818
rect 4330 77766 4342 77818
rect 4342 77766 4356 77818
rect 4380 77766 4394 77818
rect 4394 77766 4406 77818
rect 4406 77766 4436 77818
rect 4460 77766 4470 77818
rect 4470 77766 4516 77818
rect 4220 77764 4276 77766
rect 4300 77764 4356 77766
rect 4380 77764 4436 77766
rect 4460 77764 4516 77766
rect 34940 77818 34996 77820
rect 35020 77818 35076 77820
rect 35100 77818 35156 77820
rect 35180 77818 35236 77820
rect 34940 77766 34986 77818
rect 34986 77766 34996 77818
rect 35020 77766 35050 77818
rect 35050 77766 35062 77818
rect 35062 77766 35076 77818
rect 35100 77766 35114 77818
rect 35114 77766 35126 77818
rect 35126 77766 35156 77818
rect 35180 77766 35190 77818
rect 35190 77766 35236 77818
rect 34940 77764 34996 77766
rect 35020 77764 35076 77766
rect 35100 77764 35156 77766
rect 35180 77764 35236 77766
rect 4880 77274 4936 77276
rect 4960 77274 5016 77276
rect 5040 77274 5096 77276
rect 5120 77274 5176 77276
rect 4880 77222 4926 77274
rect 4926 77222 4936 77274
rect 4960 77222 4990 77274
rect 4990 77222 5002 77274
rect 5002 77222 5016 77274
rect 5040 77222 5054 77274
rect 5054 77222 5066 77274
rect 5066 77222 5096 77274
rect 5120 77222 5130 77274
rect 5130 77222 5176 77274
rect 4880 77220 4936 77222
rect 4960 77220 5016 77222
rect 5040 77220 5096 77222
rect 5120 77220 5176 77222
rect 35600 77274 35656 77276
rect 35680 77274 35736 77276
rect 35760 77274 35816 77276
rect 35840 77274 35896 77276
rect 35600 77222 35646 77274
rect 35646 77222 35656 77274
rect 35680 77222 35710 77274
rect 35710 77222 35722 77274
rect 35722 77222 35736 77274
rect 35760 77222 35774 77274
rect 35774 77222 35786 77274
rect 35786 77222 35816 77274
rect 35840 77222 35850 77274
rect 35850 77222 35896 77274
rect 35600 77220 35656 77222
rect 35680 77220 35736 77222
rect 35760 77220 35816 77222
rect 35840 77220 35896 77222
rect 4220 76730 4276 76732
rect 4300 76730 4356 76732
rect 4380 76730 4436 76732
rect 4460 76730 4516 76732
rect 4220 76678 4266 76730
rect 4266 76678 4276 76730
rect 4300 76678 4330 76730
rect 4330 76678 4342 76730
rect 4342 76678 4356 76730
rect 4380 76678 4394 76730
rect 4394 76678 4406 76730
rect 4406 76678 4436 76730
rect 4460 76678 4470 76730
rect 4470 76678 4516 76730
rect 4220 76676 4276 76678
rect 4300 76676 4356 76678
rect 4380 76676 4436 76678
rect 4460 76676 4516 76678
rect 34940 76730 34996 76732
rect 35020 76730 35076 76732
rect 35100 76730 35156 76732
rect 35180 76730 35236 76732
rect 34940 76678 34986 76730
rect 34986 76678 34996 76730
rect 35020 76678 35050 76730
rect 35050 76678 35062 76730
rect 35062 76678 35076 76730
rect 35100 76678 35114 76730
rect 35114 76678 35126 76730
rect 35126 76678 35156 76730
rect 35180 76678 35190 76730
rect 35190 76678 35236 76730
rect 34940 76676 34996 76678
rect 35020 76676 35076 76678
rect 35100 76676 35156 76678
rect 35180 76676 35236 76678
rect 4880 76186 4936 76188
rect 4960 76186 5016 76188
rect 5040 76186 5096 76188
rect 5120 76186 5176 76188
rect 4880 76134 4926 76186
rect 4926 76134 4936 76186
rect 4960 76134 4990 76186
rect 4990 76134 5002 76186
rect 5002 76134 5016 76186
rect 5040 76134 5054 76186
rect 5054 76134 5066 76186
rect 5066 76134 5096 76186
rect 5120 76134 5130 76186
rect 5130 76134 5176 76186
rect 4880 76132 4936 76134
rect 4960 76132 5016 76134
rect 5040 76132 5096 76134
rect 5120 76132 5176 76134
rect 35600 76186 35656 76188
rect 35680 76186 35736 76188
rect 35760 76186 35816 76188
rect 35840 76186 35896 76188
rect 35600 76134 35646 76186
rect 35646 76134 35656 76186
rect 35680 76134 35710 76186
rect 35710 76134 35722 76186
rect 35722 76134 35736 76186
rect 35760 76134 35774 76186
rect 35774 76134 35786 76186
rect 35786 76134 35816 76186
rect 35840 76134 35850 76186
rect 35850 76134 35896 76186
rect 35600 76132 35656 76134
rect 35680 76132 35736 76134
rect 35760 76132 35816 76134
rect 35840 76132 35896 76134
rect 4220 75642 4276 75644
rect 4300 75642 4356 75644
rect 4380 75642 4436 75644
rect 4460 75642 4516 75644
rect 4220 75590 4266 75642
rect 4266 75590 4276 75642
rect 4300 75590 4330 75642
rect 4330 75590 4342 75642
rect 4342 75590 4356 75642
rect 4380 75590 4394 75642
rect 4394 75590 4406 75642
rect 4406 75590 4436 75642
rect 4460 75590 4470 75642
rect 4470 75590 4516 75642
rect 4220 75588 4276 75590
rect 4300 75588 4356 75590
rect 4380 75588 4436 75590
rect 4460 75588 4516 75590
rect 34940 75642 34996 75644
rect 35020 75642 35076 75644
rect 35100 75642 35156 75644
rect 35180 75642 35236 75644
rect 34940 75590 34986 75642
rect 34986 75590 34996 75642
rect 35020 75590 35050 75642
rect 35050 75590 35062 75642
rect 35062 75590 35076 75642
rect 35100 75590 35114 75642
rect 35114 75590 35126 75642
rect 35126 75590 35156 75642
rect 35180 75590 35190 75642
rect 35190 75590 35236 75642
rect 34940 75588 34996 75590
rect 35020 75588 35076 75590
rect 35100 75588 35156 75590
rect 35180 75588 35236 75590
rect 4880 75098 4936 75100
rect 4960 75098 5016 75100
rect 5040 75098 5096 75100
rect 5120 75098 5176 75100
rect 4880 75046 4926 75098
rect 4926 75046 4936 75098
rect 4960 75046 4990 75098
rect 4990 75046 5002 75098
rect 5002 75046 5016 75098
rect 5040 75046 5054 75098
rect 5054 75046 5066 75098
rect 5066 75046 5096 75098
rect 5120 75046 5130 75098
rect 5130 75046 5176 75098
rect 4880 75044 4936 75046
rect 4960 75044 5016 75046
rect 5040 75044 5096 75046
rect 5120 75044 5176 75046
rect 35600 75098 35656 75100
rect 35680 75098 35736 75100
rect 35760 75098 35816 75100
rect 35840 75098 35896 75100
rect 35600 75046 35646 75098
rect 35646 75046 35656 75098
rect 35680 75046 35710 75098
rect 35710 75046 35722 75098
rect 35722 75046 35736 75098
rect 35760 75046 35774 75098
rect 35774 75046 35786 75098
rect 35786 75046 35816 75098
rect 35840 75046 35850 75098
rect 35850 75046 35896 75098
rect 35600 75044 35656 75046
rect 35680 75044 35736 75046
rect 35760 75044 35816 75046
rect 35840 75044 35896 75046
rect 4220 74554 4276 74556
rect 4300 74554 4356 74556
rect 4380 74554 4436 74556
rect 4460 74554 4516 74556
rect 4220 74502 4266 74554
rect 4266 74502 4276 74554
rect 4300 74502 4330 74554
rect 4330 74502 4342 74554
rect 4342 74502 4356 74554
rect 4380 74502 4394 74554
rect 4394 74502 4406 74554
rect 4406 74502 4436 74554
rect 4460 74502 4470 74554
rect 4470 74502 4516 74554
rect 4220 74500 4276 74502
rect 4300 74500 4356 74502
rect 4380 74500 4436 74502
rect 4460 74500 4516 74502
rect 34940 74554 34996 74556
rect 35020 74554 35076 74556
rect 35100 74554 35156 74556
rect 35180 74554 35236 74556
rect 34940 74502 34986 74554
rect 34986 74502 34996 74554
rect 35020 74502 35050 74554
rect 35050 74502 35062 74554
rect 35062 74502 35076 74554
rect 35100 74502 35114 74554
rect 35114 74502 35126 74554
rect 35126 74502 35156 74554
rect 35180 74502 35190 74554
rect 35190 74502 35236 74554
rect 34940 74500 34996 74502
rect 35020 74500 35076 74502
rect 35100 74500 35156 74502
rect 35180 74500 35236 74502
rect 4880 74010 4936 74012
rect 4960 74010 5016 74012
rect 5040 74010 5096 74012
rect 5120 74010 5176 74012
rect 4880 73958 4926 74010
rect 4926 73958 4936 74010
rect 4960 73958 4990 74010
rect 4990 73958 5002 74010
rect 5002 73958 5016 74010
rect 5040 73958 5054 74010
rect 5054 73958 5066 74010
rect 5066 73958 5096 74010
rect 5120 73958 5130 74010
rect 5130 73958 5176 74010
rect 4880 73956 4936 73958
rect 4960 73956 5016 73958
rect 5040 73956 5096 73958
rect 5120 73956 5176 73958
rect 35600 74010 35656 74012
rect 35680 74010 35736 74012
rect 35760 74010 35816 74012
rect 35840 74010 35896 74012
rect 35600 73958 35646 74010
rect 35646 73958 35656 74010
rect 35680 73958 35710 74010
rect 35710 73958 35722 74010
rect 35722 73958 35736 74010
rect 35760 73958 35774 74010
rect 35774 73958 35786 74010
rect 35786 73958 35816 74010
rect 35840 73958 35850 74010
rect 35850 73958 35896 74010
rect 35600 73956 35656 73958
rect 35680 73956 35736 73958
rect 35760 73956 35816 73958
rect 35840 73956 35896 73958
rect 4220 73466 4276 73468
rect 4300 73466 4356 73468
rect 4380 73466 4436 73468
rect 4460 73466 4516 73468
rect 4220 73414 4266 73466
rect 4266 73414 4276 73466
rect 4300 73414 4330 73466
rect 4330 73414 4342 73466
rect 4342 73414 4356 73466
rect 4380 73414 4394 73466
rect 4394 73414 4406 73466
rect 4406 73414 4436 73466
rect 4460 73414 4470 73466
rect 4470 73414 4516 73466
rect 4220 73412 4276 73414
rect 4300 73412 4356 73414
rect 4380 73412 4436 73414
rect 4460 73412 4516 73414
rect 34940 73466 34996 73468
rect 35020 73466 35076 73468
rect 35100 73466 35156 73468
rect 35180 73466 35236 73468
rect 34940 73414 34986 73466
rect 34986 73414 34996 73466
rect 35020 73414 35050 73466
rect 35050 73414 35062 73466
rect 35062 73414 35076 73466
rect 35100 73414 35114 73466
rect 35114 73414 35126 73466
rect 35126 73414 35156 73466
rect 35180 73414 35190 73466
rect 35190 73414 35236 73466
rect 34940 73412 34996 73414
rect 35020 73412 35076 73414
rect 35100 73412 35156 73414
rect 35180 73412 35236 73414
rect 4880 72922 4936 72924
rect 4960 72922 5016 72924
rect 5040 72922 5096 72924
rect 5120 72922 5176 72924
rect 4880 72870 4926 72922
rect 4926 72870 4936 72922
rect 4960 72870 4990 72922
rect 4990 72870 5002 72922
rect 5002 72870 5016 72922
rect 5040 72870 5054 72922
rect 5054 72870 5066 72922
rect 5066 72870 5096 72922
rect 5120 72870 5130 72922
rect 5130 72870 5176 72922
rect 4880 72868 4936 72870
rect 4960 72868 5016 72870
rect 5040 72868 5096 72870
rect 5120 72868 5176 72870
rect 35600 72922 35656 72924
rect 35680 72922 35736 72924
rect 35760 72922 35816 72924
rect 35840 72922 35896 72924
rect 35600 72870 35646 72922
rect 35646 72870 35656 72922
rect 35680 72870 35710 72922
rect 35710 72870 35722 72922
rect 35722 72870 35736 72922
rect 35760 72870 35774 72922
rect 35774 72870 35786 72922
rect 35786 72870 35816 72922
rect 35840 72870 35850 72922
rect 35850 72870 35896 72922
rect 35600 72868 35656 72870
rect 35680 72868 35736 72870
rect 35760 72868 35816 72870
rect 35840 72868 35896 72870
rect 4220 72378 4276 72380
rect 4300 72378 4356 72380
rect 4380 72378 4436 72380
rect 4460 72378 4516 72380
rect 4220 72326 4266 72378
rect 4266 72326 4276 72378
rect 4300 72326 4330 72378
rect 4330 72326 4342 72378
rect 4342 72326 4356 72378
rect 4380 72326 4394 72378
rect 4394 72326 4406 72378
rect 4406 72326 4436 72378
rect 4460 72326 4470 72378
rect 4470 72326 4516 72378
rect 4220 72324 4276 72326
rect 4300 72324 4356 72326
rect 4380 72324 4436 72326
rect 4460 72324 4516 72326
rect 34940 72378 34996 72380
rect 35020 72378 35076 72380
rect 35100 72378 35156 72380
rect 35180 72378 35236 72380
rect 34940 72326 34986 72378
rect 34986 72326 34996 72378
rect 35020 72326 35050 72378
rect 35050 72326 35062 72378
rect 35062 72326 35076 72378
rect 35100 72326 35114 72378
rect 35114 72326 35126 72378
rect 35126 72326 35156 72378
rect 35180 72326 35190 72378
rect 35190 72326 35236 72378
rect 34940 72324 34996 72326
rect 35020 72324 35076 72326
rect 35100 72324 35156 72326
rect 35180 72324 35236 72326
rect 4880 71834 4936 71836
rect 4960 71834 5016 71836
rect 5040 71834 5096 71836
rect 5120 71834 5176 71836
rect 4880 71782 4926 71834
rect 4926 71782 4936 71834
rect 4960 71782 4990 71834
rect 4990 71782 5002 71834
rect 5002 71782 5016 71834
rect 5040 71782 5054 71834
rect 5054 71782 5066 71834
rect 5066 71782 5096 71834
rect 5120 71782 5130 71834
rect 5130 71782 5176 71834
rect 4880 71780 4936 71782
rect 4960 71780 5016 71782
rect 5040 71780 5096 71782
rect 5120 71780 5176 71782
rect 35600 71834 35656 71836
rect 35680 71834 35736 71836
rect 35760 71834 35816 71836
rect 35840 71834 35896 71836
rect 35600 71782 35646 71834
rect 35646 71782 35656 71834
rect 35680 71782 35710 71834
rect 35710 71782 35722 71834
rect 35722 71782 35736 71834
rect 35760 71782 35774 71834
rect 35774 71782 35786 71834
rect 35786 71782 35816 71834
rect 35840 71782 35850 71834
rect 35850 71782 35896 71834
rect 35600 71780 35656 71782
rect 35680 71780 35736 71782
rect 35760 71780 35816 71782
rect 35840 71780 35896 71782
rect 4220 71290 4276 71292
rect 4300 71290 4356 71292
rect 4380 71290 4436 71292
rect 4460 71290 4516 71292
rect 4220 71238 4266 71290
rect 4266 71238 4276 71290
rect 4300 71238 4330 71290
rect 4330 71238 4342 71290
rect 4342 71238 4356 71290
rect 4380 71238 4394 71290
rect 4394 71238 4406 71290
rect 4406 71238 4436 71290
rect 4460 71238 4470 71290
rect 4470 71238 4516 71290
rect 4220 71236 4276 71238
rect 4300 71236 4356 71238
rect 4380 71236 4436 71238
rect 4460 71236 4516 71238
rect 34940 71290 34996 71292
rect 35020 71290 35076 71292
rect 35100 71290 35156 71292
rect 35180 71290 35236 71292
rect 34940 71238 34986 71290
rect 34986 71238 34996 71290
rect 35020 71238 35050 71290
rect 35050 71238 35062 71290
rect 35062 71238 35076 71290
rect 35100 71238 35114 71290
rect 35114 71238 35126 71290
rect 35126 71238 35156 71290
rect 35180 71238 35190 71290
rect 35190 71238 35236 71290
rect 34940 71236 34996 71238
rect 35020 71236 35076 71238
rect 35100 71236 35156 71238
rect 35180 71236 35236 71238
rect 4880 70746 4936 70748
rect 4960 70746 5016 70748
rect 5040 70746 5096 70748
rect 5120 70746 5176 70748
rect 4880 70694 4926 70746
rect 4926 70694 4936 70746
rect 4960 70694 4990 70746
rect 4990 70694 5002 70746
rect 5002 70694 5016 70746
rect 5040 70694 5054 70746
rect 5054 70694 5066 70746
rect 5066 70694 5096 70746
rect 5120 70694 5130 70746
rect 5130 70694 5176 70746
rect 4880 70692 4936 70694
rect 4960 70692 5016 70694
rect 5040 70692 5096 70694
rect 5120 70692 5176 70694
rect 35600 70746 35656 70748
rect 35680 70746 35736 70748
rect 35760 70746 35816 70748
rect 35840 70746 35896 70748
rect 35600 70694 35646 70746
rect 35646 70694 35656 70746
rect 35680 70694 35710 70746
rect 35710 70694 35722 70746
rect 35722 70694 35736 70746
rect 35760 70694 35774 70746
rect 35774 70694 35786 70746
rect 35786 70694 35816 70746
rect 35840 70694 35850 70746
rect 35850 70694 35896 70746
rect 35600 70692 35656 70694
rect 35680 70692 35736 70694
rect 35760 70692 35816 70694
rect 35840 70692 35896 70694
rect 4220 70202 4276 70204
rect 4300 70202 4356 70204
rect 4380 70202 4436 70204
rect 4460 70202 4516 70204
rect 4220 70150 4266 70202
rect 4266 70150 4276 70202
rect 4300 70150 4330 70202
rect 4330 70150 4342 70202
rect 4342 70150 4356 70202
rect 4380 70150 4394 70202
rect 4394 70150 4406 70202
rect 4406 70150 4436 70202
rect 4460 70150 4470 70202
rect 4470 70150 4516 70202
rect 4220 70148 4276 70150
rect 4300 70148 4356 70150
rect 4380 70148 4436 70150
rect 4460 70148 4516 70150
rect 34940 70202 34996 70204
rect 35020 70202 35076 70204
rect 35100 70202 35156 70204
rect 35180 70202 35236 70204
rect 34940 70150 34986 70202
rect 34986 70150 34996 70202
rect 35020 70150 35050 70202
rect 35050 70150 35062 70202
rect 35062 70150 35076 70202
rect 35100 70150 35114 70202
rect 35114 70150 35126 70202
rect 35126 70150 35156 70202
rect 35180 70150 35190 70202
rect 35190 70150 35236 70202
rect 34940 70148 34996 70150
rect 35020 70148 35076 70150
rect 35100 70148 35156 70150
rect 35180 70148 35236 70150
rect 4880 69658 4936 69660
rect 4960 69658 5016 69660
rect 5040 69658 5096 69660
rect 5120 69658 5176 69660
rect 4880 69606 4926 69658
rect 4926 69606 4936 69658
rect 4960 69606 4990 69658
rect 4990 69606 5002 69658
rect 5002 69606 5016 69658
rect 5040 69606 5054 69658
rect 5054 69606 5066 69658
rect 5066 69606 5096 69658
rect 5120 69606 5130 69658
rect 5130 69606 5176 69658
rect 4880 69604 4936 69606
rect 4960 69604 5016 69606
rect 5040 69604 5096 69606
rect 5120 69604 5176 69606
rect 35600 69658 35656 69660
rect 35680 69658 35736 69660
rect 35760 69658 35816 69660
rect 35840 69658 35896 69660
rect 35600 69606 35646 69658
rect 35646 69606 35656 69658
rect 35680 69606 35710 69658
rect 35710 69606 35722 69658
rect 35722 69606 35736 69658
rect 35760 69606 35774 69658
rect 35774 69606 35786 69658
rect 35786 69606 35816 69658
rect 35840 69606 35850 69658
rect 35850 69606 35896 69658
rect 35600 69604 35656 69606
rect 35680 69604 35736 69606
rect 35760 69604 35816 69606
rect 35840 69604 35896 69606
rect 4220 69114 4276 69116
rect 4300 69114 4356 69116
rect 4380 69114 4436 69116
rect 4460 69114 4516 69116
rect 4220 69062 4266 69114
rect 4266 69062 4276 69114
rect 4300 69062 4330 69114
rect 4330 69062 4342 69114
rect 4342 69062 4356 69114
rect 4380 69062 4394 69114
rect 4394 69062 4406 69114
rect 4406 69062 4436 69114
rect 4460 69062 4470 69114
rect 4470 69062 4516 69114
rect 4220 69060 4276 69062
rect 4300 69060 4356 69062
rect 4380 69060 4436 69062
rect 4460 69060 4516 69062
rect 34940 69114 34996 69116
rect 35020 69114 35076 69116
rect 35100 69114 35156 69116
rect 35180 69114 35236 69116
rect 34940 69062 34986 69114
rect 34986 69062 34996 69114
rect 35020 69062 35050 69114
rect 35050 69062 35062 69114
rect 35062 69062 35076 69114
rect 35100 69062 35114 69114
rect 35114 69062 35126 69114
rect 35126 69062 35156 69114
rect 35180 69062 35190 69114
rect 35190 69062 35236 69114
rect 34940 69060 34996 69062
rect 35020 69060 35076 69062
rect 35100 69060 35156 69062
rect 35180 69060 35236 69062
rect 4880 68570 4936 68572
rect 4960 68570 5016 68572
rect 5040 68570 5096 68572
rect 5120 68570 5176 68572
rect 4880 68518 4926 68570
rect 4926 68518 4936 68570
rect 4960 68518 4990 68570
rect 4990 68518 5002 68570
rect 5002 68518 5016 68570
rect 5040 68518 5054 68570
rect 5054 68518 5066 68570
rect 5066 68518 5096 68570
rect 5120 68518 5130 68570
rect 5130 68518 5176 68570
rect 4880 68516 4936 68518
rect 4960 68516 5016 68518
rect 5040 68516 5096 68518
rect 5120 68516 5176 68518
rect 35600 68570 35656 68572
rect 35680 68570 35736 68572
rect 35760 68570 35816 68572
rect 35840 68570 35896 68572
rect 35600 68518 35646 68570
rect 35646 68518 35656 68570
rect 35680 68518 35710 68570
rect 35710 68518 35722 68570
rect 35722 68518 35736 68570
rect 35760 68518 35774 68570
rect 35774 68518 35786 68570
rect 35786 68518 35816 68570
rect 35840 68518 35850 68570
rect 35850 68518 35896 68570
rect 35600 68516 35656 68518
rect 35680 68516 35736 68518
rect 35760 68516 35816 68518
rect 35840 68516 35896 68518
rect 4220 68026 4276 68028
rect 4300 68026 4356 68028
rect 4380 68026 4436 68028
rect 4460 68026 4516 68028
rect 4220 67974 4266 68026
rect 4266 67974 4276 68026
rect 4300 67974 4330 68026
rect 4330 67974 4342 68026
rect 4342 67974 4356 68026
rect 4380 67974 4394 68026
rect 4394 67974 4406 68026
rect 4406 67974 4436 68026
rect 4460 67974 4470 68026
rect 4470 67974 4516 68026
rect 4220 67972 4276 67974
rect 4300 67972 4356 67974
rect 4380 67972 4436 67974
rect 4460 67972 4516 67974
rect 34940 68026 34996 68028
rect 35020 68026 35076 68028
rect 35100 68026 35156 68028
rect 35180 68026 35236 68028
rect 34940 67974 34986 68026
rect 34986 67974 34996 68026
rect 35020 67974 35050 68026
rect 35050 67974 35062 68026
rect 35062 67974 35076 68026
rect 35100 67974 35114 68026
rect 35114 67974 35126 68026
rect 35126 67974 35156 68026
rect 35180 67974 35190 68026
rect 35190 67974 35236 68026
rect 34940 67972 34996 67974
rect 35020 67972 35076 67974
rect 35100 67972 35156 67974
rect 35180 67972 35236 67974
rect 4880 67482 4936 67484
rect 4960 67482 5016 67484
rect 5040 67482 5096 67484
rect 5120 67482 5176 67484
rect 4880 67430 4926 67482
rect 4926 67430 4936 67482
rect 4960 67430 4990 67482
rect 4990 67430 5002 67482
rect 5002 67430 5016 67482
rect 5040 67430 5054 67482
rect 5054 67430 5066 67482
rect 5066 67430 5096 67482
rect 5120 67430 5130 67482
rect 5130 67430 5176 67482
rect 4880 67428 4936 67430
rect 4960 67428 5016 67430
rect 5040 67428 5096 67430
rect 5120 67428 5176 67430
rect 35600 67482 35656 67484
rect 35680 67482 35736 67484
rect 35760 67482 35816 67484
rect 35840 67482 35896 67484
rect 35600 67430 35646 67482
rect 35646 67430 35656 67482
rect 35680 67430 35710 67482
rect 35710 67430 35722 67482
rect 35722 67430 35736 67482
rect 35760 67430 35774 67482
rect 35774 67430 35786 67482
rect 35786 67430 35816 67482
rect 35840 67430 35850 67482
rect 35850 67430 35896 67482
rect 35600 67428 35656 67430
rect 35680 67428 35736 67430
rect 35760 67428 35816 67430
rect 35840 67428 35896 67430
rect 4220 66938 4276 66940
rect 4300 66938 4356 66940
rect 4380 66938 4436 66940
rect 4460 66938 4516 66940
rect 4220 66886 4266 66938
rect 4266 66886 4276 66938
rect 4300 66886 4330 66938
rect 4330 66886 4342 66938
rect 4342 66886 4356 66938
rect 4380 66886 4394 66938
rect 4394 66886 4406 66938
rect 4406 66886 4436 66938
rect 4460 66886 4470 66938
rect 4470 66886 4516 66938
rect 4220 66884 4276 66886
rect 4300 66884 4356 66886
rect 4380 66884 4436 66886
rect 4460 66884 4516 66886
rect 34940 66938 34996 66940
rect 35020 66938 35076 66940
rect 35100 66938 35156 66940
rect 35180 66938 35236 66940
rect 34940 66886 34986 66938
rect 34986 66886 34996 66938
rect 35020 66886 35050 66938
rect 35050 66886 35062 66938
rect 35062 66886 35076 66938
rect 35100 66886 35114 66938
rect 35114 66886 35126 66938
rect 35126 66886 35156 66938
rect 35180 66886 35190 66938
rect 35190 66886 35236 66938
rect 34940 66884 34996 66886
rect 35020 66884 35076 66886
rect 35100 66884 35156 66886
rect 35180 66884 35236 66886
rect 4880 66394 4936 66396
rect 4960 66394 5016 66396
rect 5040 66394 5096 66396
rect 5120 66394 5176 66396
rect 4880 66342 4926 66394
rect 4926 66342 4936 66394
rect 4960 66342 4990 66394
rect 4990 66342 5002 66394
rect 5002 66342 5016 66394
rect 5040 66342 5054 66394
rect 5054 66342 5066 66394
rect 5066 66342 5096 66394
rect 5120 66342 5130 66394
rect 5130 66342 5176 66394
rect 4880 66340 4936 66342
rect 4960 66340 5016 66342
rect 5040 66340 5096 66342
rect 5120 66340 5176 66342
rect 35600 66394 35656 66396
rect 35680 66394 35736 66396
rect 35760 66394 35816 66396
rect 35840 66394 35896 66396
rect 35600 66342 35646 66394
rect 35646 66342 35656 66394
rect 35680 66342 35710 66394
rect 35710 66342 35722 66394
rect 35722 66342 35736 66394
rect 35760 66342 35774 66394
rect 35774 66342 35786 66394
rect 35786 66342 35816 66394
rect 35840 66342 35850 66394
rect 35850 66342 35896 66394
rect 35600 66340 35656 66342
rect 35680 66340 35736 66342
rect 35760 66340 35816 66342
rect 35840 66340 35896 66342
rect 4220 65850 4276 65852
rect 4300 65850 4356 65852
rect 4380 65850 4436 65852
rect 4460 65850 4516 65852
rect 4220 65798 4266 65850
rect 4266 65798 4276 65850
rect 4300 65798 4330 65850
rect 4330 65798 4342 65850
rect 4342 65798 4356 65850
rect 4380 65798 4394 65850
rect 4394 65798 4406 65850
rect 4406 65798 4436 65850
rect 4460 65798 4470 65850
rect 4470 65798 4516 65850
rect 4220 65796 4276 65798
rect 4300 65796 4356 65798
rect 4380 65796 4436 65798
rect 4460 65796 4516 65798
rect 34940 65850 34996 65852
rect 35020 65850 35076 65852
rect 35100 65850 35156 65852
rect 35180 65850 35236 65852
rect 34940 65798 34986 65850
rect 34986 65798 34996 65850
rect 35020 65798 35050 65850
rect 35050 65798 35062 65850
rect 35062 65798 35076 65850
rect 35100 65798 35114 65850
rect 35114 65798 35126 65850
rect 35126 65798 35156 65850
rect 35180 65798 35190 65850
rect 35190 65798 35236 65850
rect 34940 65796 34996 65798
rect 35020 65796 35076 65798
rect 35100 65796 35156 65798
rect 35180 65796 35236 65798
rect 4880 65306 4936 65308
rect 4960 65306 5016 65308
rect 5040 65306 5096 65308
rect 5120 65306 5176 65308
rect 4880 65254 4926 65306
rect 4926 65254 4936 65306
rect 4960 65254 4990 65306
rect 4990 65254 5002 65306
rect 5002 65254 5016 65306
rect 5040 65254 5054 65306
rect 5054 65254 5066 65306
rect 5066 65254 5096 65306
rect 5120 65254 5130 65306
rect 5130 65254 5176 65306
rect 4880 65252 4936 65254
rect 4960 65252 5016 65254
rect 5040 65252 5096 65254
rect 5120 65252 5176 65254
rect 35600 65306 35656 65308
rect 35680 65306 35736 65308
rect 35760 65306 35816 65308
rect 35840 65306 35896 65308
rect 35600 65254 35646 65306
rect 35646 65254 35656 65306
rect 35680 65254 35710 65306
rect 35710 65254 35722 65306
rect 35722 65254 35736 65306
rect 35760 65254 35774 65306
rect 35774 65254 35786 65306
rect 35786 65254 35816 65306
rect 35840 65254 35850 65306
rect 35850 65254 35896 65306
rect 35600 65252 35656 65254
rect 35680 65252 35736 65254
rect 35760 65252 35816 65254
rect 35840 65252 35896 65254
rect 4220 64762 4276 64764
rect 4300 64762 4356 64764
rect 4380 64762 4436 64764
rect 4460 64762 4516 64764
rect 4220 64710 4266 64762
rect 4266 64710 4276 64762
rect 4300 64710 4330 64762
rect 4330 64710 4342 64762
rect 4342 64710 4356 64762
rect 4380 64710 4394 64762
rect 4394 64710 4406 64762
rect 4406 64710 4436 64762
rect 4460 64710 4470 64762
rect 4470 64710 4516 64762
rect 4220 64708 4276 64710
rect 4300 64708 4356 64710
rect 4380 64708 4436 64710
rect 4460 64708 4516 64710
rect 34940 64762 34996 64764
rect 35020 64762 35076 64764
rect 35100 64762 35156 64764
rect 35180 64762 35236 64764
rect 34940 64710 34986 64762
rect 34986 64710 34996 64762
rect 35020 64710 35050 64762
rect 35050 64710 35062 64762
rect 35062 64710 35076 64762
rect 35100 64710 35114 64762
rect 35114 64710 35126 64762
rect 35126 64710 35156 64762
rect 35180 64710 35190 64762
rect 35190 64710 35236 64762
rect 34940 64708 34996 64710
rect 35020 64708 35076 64710
rect 35100 64708 35156 64710
rect 35180 64708 35236 64710
rect 4880 64218 4936 64220
rect 4960 64218 5016 64220
rect 5040 64218 5096 64220
rect 5120 64218 5176 64220
rect 4880 64166 4926 64218
rect 4926 64166 4936 64218
rect 4960 64166 4990 64218
rect 4990 64166 5002 64218
rect 5002 64166 5016 64218
rect 5040 64166 5054 64218
rect 5054 64166 5066 64218
rect 5066 64166 5096 64218
rect 5120 64166 5130 64218
rect 5130 64166 5176 64218
rect 4880 64164 4936 64166
rect 4960 64164 5016 64166
rect 5040 64164 5096 64166
rect 5120 64164 5176 64166
rect 35600 64218 35656 64220
rect 35680 64218 35736 64220
rect 35760 64218 35816 64220
rect 35840 64218 35896 64220
rect 35600 64166 35646 64218
rect 35646 64166 35656 64218
rect 35680 64166 35710 64218
rect 35710 64166 35722 64218
rect 35722 64166 35736 64218
rect 35760 64166 35774 64218
rect 35774 64166 35786 64218
rect 35786 64166 35816 64218
rect 35840 64166 35850 64218
rect 35850 64166 35896 64218
rect 35600 64164 35656 64166
rect 35680 64164 35736 64166
rect 35760 64164 35816 64166
rect 35840 64164 35896 64166
rect 4220 63674 4276 63676
rect 4300 63674 4356 63676
rect 4380 63674 4436 63676
rect 4460 63674 4516 63676
rect 4220 63622 4266 63674
rect 4266 63622 4276 63674
rect 4300 63622 4330 63674
rect 4330 63622 4342 63674
rect 4342 63622 4356 63674
rect 4380 63622 4394 63674
rect 4394 63622 4406 63674
rect 4406 63622 4436 63674
rect 4460 63622 4470 63674
rect 4470 63622 4516 63674
rect 4220 63620 4276 63622
rect 4300 63620 4356 63622
rect 4380 63620 4436 63622
rect 4460 63620 4516 63622
rect 34940 63674 34996 63676
rect 35020 63674 35076 63676
rect 35100 63674 35156 63676
rect 35180 63674 35236 63676
rect 34940 63622 34986 63674
rect 34986 63622 34996 63674
rect 35020 63622 35050 63674
rect 35050 63622 35062 63674
rect 35062 63622 35076 63674
rect 35100 63622 35114 63674
rect 35114 63622 35126 63674
rect 35126 63622 35156 63674
rect 35180 63622 35190 63674
rect 35190 63622 35236 63674
rect 34940 63620 34996 63622
rect 35020 63620 35076 63622
rect 35100 63620 35156 63622
rect 35180 63620 35236 63622
rect 4880 63130 4936 63132
rect 4960 63130 5016 63132
rect 5040 63130 5096 63132
rect 5120 63130 5176 63132
rect 4880 63078 4926 63130
rect 4926 63078 4936 63130
rect 4960 63078 4990 63130
rect 4990 63078 5002 63130
rect 5002 63078 5016 63130
rect 5040 63078 5054 63130
rect 5054 63078 5066 63130
rect 5066 63078 5096 63130
rect 5120 63078 5130 63130
rect 5130 63078 5176 63130
rect 4880 63076 4936 63078
rect 4960 63076 5016 63078
rect 5040 63076 5096 63078
rect 5120 63076 5176 63078
rect 35600 63130 35656 63132
rect 35680 63130 35736 63132
rect 35760 63130 35816 63132
rect 35840 63130 35896 63132
rect 35600 63078 35646 63130
rect 35646 63078 35656 63130
rect 35680 63078 35710 63130
rect 35710 63078 35722 63130
rect 35722 63078 35736 63130
rect 35760 63078 35774 63130
rect 35774 63078 35786 63130
rect 35786 63078 35816 63130
rect 35840 63078 35850 63130
rect 35850 63078 35896 63130
rect 35600 63076 35656 63078
rect 35680 63076 35736 63078
rect 35760 63076 35816 63078
rect 35840 63076 35896 63078
rect 43626 76236 43628 76256
rect 43628 76236 43680 76256
rect 43680 76236 43682 76256
rect 43626 76200 43682 76236
rect 47950 75928 48006 75984
rect 49606 77052 49608 77072
rect 49608 77052 49660 77072
rect 49660 77052 49662 77072
rect 49606 77016 49662 77052
rect 45742 74568 45798 74624
rect 41786 62736 41842 62792
rect 4220 62586 4276 62588
rect 4300 62586 4356 62588
rect 4380 62586 4436 62588
rect 4460 62586 4516 62588
rect 4220 62534 4266 62586
rect 4266 62534 4276 62586
rect 4300 62534 4330 62586
rect 4330 62534 4342 62586
rect 4342 62534 4356 62586
rect 4380 62534 4394 62586
rect 4394 62534 4406 62586
rect 4406 62534 4436 62586
rect 4460 62534 4470 62586
rect 4470 62534 4516 62586
rect 4220 62532 4276 62534
rect 4300 62532 4356 62534
rect 4380 62532 4436 62534
rect 4460 62532 4516 62534
rect 34940 62586 34996 62588
rect 35020 62586 35076 62588
rect 35100 62586 35156 62588
rect 35180 62586 35236 62588
rect 34940 62534 34986 62586
rect 34986 62534 34996 62586
rect 35020 62534 35050 62586
rect 35050 62534 35062 62586
rect 35062 62534 35076 62586
rect 35100 62534 35114 62586
rect 35114 62534 35126 62586
rect 35126 62534 35156 62586
rect 35180 62534 35190 62586
rect 35190 62534 35236 62586
rect 34940 62532 34996 62534
rect 35020 62532 35076 62534
rect 35100 62532 35156 62534
rect 35180 62532 35236 62534
rect 1490 61920 1546 61976
rect 846 61376 902 61432
rect 4880 62042 4936 62044
rect 4960 62042 5016 62044
rect 5040 62042 5096 62044
rect 5120 62042 5176 62044
rect 4880 61990 4926 62042
rect 4926 61990 4936 62042
rect 4960 61990 4990 62042
rect 4990 61990 5002 62042
rect 5002 61990 5016 62042
rect 5040 61990 5054 62042
rect 5054 61990 5066 62042
rect 5066 61990 5096 62042
rect 5120 61990 5130 62042
rect 5130 61990 5176 62042
rect 4880 61988 4936 61990
rect 4960 61988 5016 61990
rect 5040 61988 5096 61990
rect 5120 61988 5176 61990
rect 35600 62042 35656 62044
rect 35680 62042 35736 62044
rect 35760 62042 35816 62044
rect 35840 62042 35896 62044
rect 35600 61990 35646 62042
rect 35646 61990 35656 62042
rect 35680 61990 35710 62042
rect 35710 61990 35722 62042
rect 35722 61990 35736 62042
rect 35760 61990 35774 62042
rect 35774 61990 35786 62042
rect 35786 61990 35816 62042
rect 35840 61990 35850 62042
rect 35850 61990 35896 62042
rect 35600 61988 35656 61990
rect 35680 61988 35736 61990
rect 35760 61988 35816 61990
rect 35840 61988 35896 61990
rect 4220 61498 4276 61500
rect 4300 61498 4356 61500
rect 4380 61498 4436 61500
rect 4460 61498 4516 61500
rect 4220 61446 4266 61498
rect 4266 61446 4276 61498
rect 4300 61446 4330 61498
rect 4330 61446 4342 61498
rect 4342 61446 4356 61498
rect 4380 61446 4394 61498
rect 4394 61446 4406 61498
rect 4406 61446 4436 61498
rect 4460 61446 4470 61498
rect 4470 61446 4516 61498
rect 4220 61444 4276 61446
rect 4300 61444 4356 61446
rect 4380 61444 4436 61446
rect 4460 61444 4516 61446
rect 34940 61498 34996 61500
rect 35020 61498 35076 61500
rect 35100 61498 35156 61500
rect 35180 61498 35236 61500
rect 34940 61446 34986 61498
rect 34986 61446 34996 61498
rect 35020 61446 35050 61498
rect 35050 61446 35062 61498
rect 35062 61446 35076 61498
rect 35100 61446 35114 61498
rect 35114 61446 35126 61498
rect 35126 61446 35156 61498
rect 35180 61446 35190 61498
rect 35190 61446 35236 61498
rect 34940 61444 34996 61446
rect 35020 61444 35076 61446
rect 35100 61444 35156 61446
rect 35180 61444 35236 61446
rect 4880 60954 4936 60956
rect 4960 60954 5016 60956
rect 5040 60954 5096 60956
rect 5120 60954 5176 60956
rect 4880 60902 4926 60954
rect 4926 60902 4936 60954
rect 4960 60902 4990 60954
rect 4990 60902 5002 60954
rect 5002 60902 5016 60954
rect 5040 60902 5054 60954
rect 5054 60902 5066 60954
rect 5066 60902 5096 60954
rect 5120 60902 5130 60954
rect 5130 60902 5176 60954
rect 4880 60900 4936 60902
rect 4960 60900 5016 60902
rect 5040 60900 5096 60902
rect 5120 60900 5176 60902
rect 1312 60410 1368 60412
rect 1392 60410 1448 60412
rect 1312 60358 1322 60410
rect 1322 60358 1368 60410
rect 1392 60358 1438 60410
rect 1438 60358 1448 60410
rect 1312 60356 1368 60358
rect 1392 60356 1448 60358
rect 4220 60410 4276 60412
rect 4300 60410 4356 60412
rect 4380 60410 4436 60412
rect 4460 60410 4516 60412
rect 4220 60358 4266 60410
rect 4266 60358 4276 60410
rect 4300 60358 4330 60410
rect 4330 60358 4342 60410
rect 4342 60358 4356 60410
rect 4380 60358 4394 60410
rect 4394 60358 4406 60410
rect 4406 60358 4436 60410
rect 4460 60358 4470 60410
rect 4470 60358 4516 60410
rect 4220 60356 4276 60358
rect 4300 60356 4356 60358
rect 4380 60356 4436 60358
rect 4460 60356 4516 60358
rect 1680 59866 1736 59868
rect 1760 59866 1816 59868
rect 1680 59814 1690 59866
rect 1690 59814 1736 59866
rect 1760 59814 1806 59866
rect 1806 59814 1816 59866
rect 1680 59812 1736 59814
rect 1760 59812 1816 59814
rect 4880 59866 4936 59868
rect 4960 59866 5016 59868
rect 5040 59866 5096 59868
rect 5120 59866 5176 59868
rect 4880 59814 4926 59866
rect 4926 59814 4936 59866
rect 4960 59814 4990 59866
rect 4990 59814 5002 59866
rect 5002 59814 5016 59866
rect 5040 59814 5054 59866
rect 5054 59814 5066 59866
rect 5066 59814 5096 59866
rect 5120 59814 5130 59866
rect 5130 59814 5176 59866
rect 4880 59812 4936 59814
rect 4960 59812 5016 59814
rect 5040 59812 5096 59814
rect 5120 59812 5176 59814
rect 1312 59322 1368 59324
rect 1392 59322 1448 59324
rect 1312 59270 1322 59322
rect 1322 59270 1368 59322
rect 1392 59270 1438 59322
rect 1438 59270 1448 59322
rect 1312 59268 1368 59270
rect 1392 59268 1448 59270
rect 1680 58778 1736 58780
rect 1760 58778 1816 58780
rect 1680 58726 1690 58778
rect 1690 58726 1736 58778
rect 1760 58726 1806 58778
rect 1806 58726 1816 58778
rect 1680 58724 1736 58726
rect 1760 58724 1816 58726
rect 1312 58234 1368 58236
rect 1392 58234 1448 58236
rect 1312 58182 1322 58234
rect 1322 58182 1368 58234
rect 1392 58182 1438 58234
rect 1438 58182 1448 58234
rect 1312 58180 1368 58182
rect 1392 58180 1448 58182
rect 1680 57690 1736 57692
rect 1760 57690 1816 57692
rect 1680 57638 1690 57690
rect 1690 57638 1736 57690
rect 1760 57638 1806 57690
rect 1806 57638 1816 57690
rect 1680 57636 1736 57638
rect 1760 57636 1816 57638
rect 1312 57146 1368 57148
rect 1392 57146 1448 57148
rect 1312 57094 1322 57146
rect 1322 57094 1368 57146
rect 1392 57094 1438 57146
rect 1438 57094 1448 57146
rect 1312 57092 1368 57094
rect 1392 57092 1448 57094
rect 1680 56602 1736 56604
rect 1760 56602 1816 56604
rect 1680 56550 1690 56602
rect 1690 56550 1736 56602
rect 1760 56550 1806 56602
rect 1806 56550 1816 56602
rect 1680 56548 1736 56550
rect 1760 56548 1816 56550
rect 1312 56058 1368 56060
rect 1392 56058 1448 56060
rect 1312 56006 1322 56058
rect 1322 56006 1368 56058
rect 1392 56006 1438 56058
rect 1438 56006 1448 56058
rect 1312 56004 1368 56006
rect 1392 56004 1448 56006
rect 1680 55514 1736 55516
rect 1760 55514 1816 55516
rect 1680 55462 1690 55514
rect 1690 55462 1736 55514
rect 1760 55462 1806 55514
rect 1806 55462 1816 55514
rect 1680 55460 1736 55462
rect 1760 55460 1816 55462
rect 1312 54970 1368 54972
rect 1392 54970 1448 54972
rect 1312 54918 1322 54970
rect 1322 54918 1368 54970
rect 1392 54918 1438 54970
rect 1438 54918 1448 54970
rect 1312 54916 1368 54918
rect 1392 54916 1448 54918
rect 1680 54426 1736 54428
rect 1760 54426 1816 54428
rect 1680 54374 1690 54426
rect 1690 54374 1736 54426
rect 1760 54374 1806 54426
rect 1806 54374 1816 54426
rect 1680 54372 1736 54374
rect 1760 54372 1816 54374
rect 1312 53882 1368 53884
rect 1392 53882 1448 53884
rect 1312 53830 1322 53882
rect 1322 53830 1368 53882
rect 1392 53830 1438 53882
rect 1438 53830 1448 53882
rect 1312 53828 1368 53830
rect 1392 53828 1448 53830
rect 1680 53338 1736 53340
rect 1760 53338 1816 53340
rect 1680 53286 1690 53338
rect 1690 53286 1736 53338
rect 1760 53286 1806 53338
rect 1806 53286 1816 53338
rect 1680 53284 1736 53286
rect 1760 53284 1816 53286
rect 1312 52794 1368 52796
rect 1392 52794 1448 52796
rect 1312 52742 1322 52794
rect 1322 52742 1368 52794
rect 1392 52742 1438 52794
rect 1438 52742 1448 52794
rect 1312 52740 1368 52742
rect 1392 52740 1448 52742
rect 1680 52250 1736 52252
rect 1760 52250 1816 52252
rect 1680 52198 1690 52250
rect 1690 52198 1736 52250
rect 1760 52198 1806 52250
rect 1806 52198 1816 52250
rect 1680 52196 1736 52198
rect 1760 52196 1816 52198
rect 1312 51706 1368 51708
rect 1392 51706 1448 51708
rect 1312 51654 1322 51706
rect 1322 51654 1368 51706
rect 1392 51654 1438 51706
rect 1438 51654 1448 51706
rect 1312 51652 1368 51654
rect 1392 51652 1448 51654
rect 1680 51162 1736 51164
rect 1760 51162 1816 51164
rect 1680 51110 1690 51162
rect 1690 51110 1736 51162
rect 1760 51110 1806 51162
rect 1806 51110 1816 51162
rect 1680 51108 1736 51110
rect 1760 51108 1816 51110
rect 1312 50618 1368 50620
rect 1392 50618 1448 50620
rect 1312 50566 1322 50618
rect 1322 50566 1368 50618
rect 1392 50566 1438 50618
rect 1438 50566 1448 50618
rect 1312 50564 1368 50566
rect 1392 50564 1448 50566
rect 1680 50074 1736 50076
rect 1760 50074 1816 50076
rect 1680 50022 1690 50074
rect 1690 50022 1736 50074
rect 1760 50022 1806 50074
rect 1806 50022 1816 50074
rect 1680 50020 1736 50022
rect 1760 50020 1816 50022
rect 1312 49530 1368 49532
rect 1392 49530 1448 49532
rect 1312 49478 1322 49530
rect 1322 49478 1368 49530
rect 1392 49478 1438 49530
rect 1438 49478 1448 49530
rect 1312 49476 1368 49478
rect 1392 49476 1448 49478
rect 1680 48986 1736 48988
rect 1760 48986 1816 48988
rect 1680 48934 1690 48986
rect 1690 48934 1736 48986
rect 1760 48934 1806 48986
rect 1806 48934 1816 48986
rect 1680 48932 1736 48934
rect 1760 48932 1816 48934
rect 1312 48442 1368 48444
rect 1392 48442 1448 48444
rect 1312 48390 1322 48442
rect 1322 48390 1368 48442
rect 1392 48390 1438 48442
rect 1438 48390 1448 48442
rect 1312 48388 1368 48390
rect 1392 48388 1448 48390
rect 1680 47898 1736 47900
rect 1760 47898 1816 47900
rect 1680 47846 1690 47898
rect 1690 47846 1736 47898
rect 1760 47846 1806 47898
rect 1806 47846 1816 47898
rect 1680 47844 1736 47846
rect 1760 47844 1816 47846
rect 1312 47354 1368 47356
rect 1392 47354 1448 47356
rect 1312 47302 1322 47354
rect 1322 47302 1368 47354
rect 1392 47302 1438 47354
rect 1438 47302 1448 47354
rect 1312 47300 1368 47302
rect 1392 47300 1448 47302
rect 1680 46810 1736 46812
rect 1760 46810 1816 46812
rect 1680 46758 1690 46810
rect 1690 46758 1736 46810
rect 1760 46758 1806 46810
rect 1806 46758 1816 46810
rect 1680 46756 1736 46758
rect 1760 46756 1816 46758
rect 1312 46266 1368 46268
rect 1392 46266 1448 46268
rect 1312 46214 1322 46266
rect 1322 46214 1368 46266
rect 1392 46214 1438 46266
rect 1438 46214 1448 46266
rect 1312 46212 1368 46214
rect 1392 46212 1448 46214
rect 1680 45722 1736 45724
rect 1760 45722 1816 45724
rect 1680 45670 1690 45722
rect 1690 45670 1736 45722
rect 1760 45670 1806 45722
rect 1806 45670 1816 45722
rect 1680 45668 1736 45670
rect 1760 45668 1816 45670
rect 1312 45178 1368 45180
rect 1392 45178 1448 45180
rect 1312 45126 1322 45178
rect 1322 45126 1368 45178
rect 1392 45126 1438 45178
rect 1438 45126 1448 45178
rect 1312 45124 1368 45126
rect 1392 45124 1448 45126
rect 1680 44634 1736 44636
rect 1760 44634 1816 44636
rect 1680 44582 1690 44634
rect 1690 44582 1736 44634
rect 1760 44582 1806 44634
rect 1806 44582 1816 44634
rect 1680 44580 1736 44582
rect 1760 44580 1816 44582
rect 1312 44090 1368 44092
rect 1392 44090 1448 44092
rect 1312 44038 1322 44090
rect 1322 44038 1368 44090
rect 1392 44038 1438 44090
rect 1438 44038 1448 44090
rect 1312 44036 1368 44038
rect 1392 44036 1448 44038
rect 1680 43546 1736 43548
rect 1760 43546 1816 43548
rect 1680 43494 1690 43546
rect 1690 43494 1736 43546
rect 1760 43494 1806 43546
rect 1806 43494 1816 43546
rect 1680 43492 1736 43494
rect 1760 43492 1816 43494
rect 1312 43002 1368 43004
rect 1392 43002 1448 43004
rect 1312 42950 1322 43002
rect 1322 42950 1368 43002
rect 1392 42950 1438 43002
rect 1438 42950 1448 43002
rect 1312 42948 1368 42950
rect 1392 42948 1448 42950
rect 1680 42458 1736 42460
rect 1760 42458 1816 42460
rect 1680 42406 1690 42458
rect 1690 42406 1736 42458
rect 1760 42406 1806 42458
rect 1806 42406 1816 42458
rect 1680 42404 1736 42406
rect 1760 42404 1816 42406
rect 1312 41914 1368 41916
rect 1392 41914 1448 41916
rect 1312 41862 1322 41914
rect 1322 41862 1368 41914
rect 1392 41862 1438 41914
rect 1438 41862 1448 41914
rect 1312 41860 1368 41862
rect 1392 41860 1448 41862
rect 1680 41370 1736 41372
rect 1760 41370 1816 41372
rect 1680 41318 1690 41370
rect 1690 41318 1736 41370
rect 1760 41318 1806 41370
rect 1806 41318 1816 41370
rect 1680 41316 1736 41318
rect 1760 41316 1816 41318
rect 1312 40826 1368 40828
rect 1392 40826 1448 40828
rect 1312 40774 1322 40826
rect 1322 40774 1368 40826
rect 1392 40774 1438 40826
rect 1438 40774 1448 40826
rect 1312 40772 1368 40774
rect 1392 40772 1448 40774
rect 1680 40282 1736 40284
rect 1760 40282 1816 40284
rect 1680 40230 1690 40282
rect 1690 40230 1736 40282
rect 1760 40230 1806 40282
rect 1806 40230 1816 40282
rect 1680 40228 1736 40230
rect 1760 40228 1816 40230
rect 1312 39738 1368 39740
rect 1392 39738 1448 39740
rect 1312 39686 1322 39738
rect 1322 39686 1368 39738
rect 1392 39686 1438 39738
rect 1438 39686 1448 39738
rect 1312 39684 1368 39686
rect 1392 39684 1448 39686
rect 1680 39194 1736 39196
rect 1760 39194 1816 39196
rect 1680 39142 1690 39194
rect 1690 39142 1736 39194
rect 1760 39142 1806 39194
rect 1806 39142 1816 39194
rect 1680 39140 1736 39142
rect 1760 39140 1816 39142
rect 1312 38650 1368 38652
rect 1392 38650 1448 38652
rect 1312 38598 1322 38650
rect 1322 38598 1368 38650
rect 1392 38598 1438 38650
rect 1438 38598 1448 38650
rect 1312 38596 1368 38598
rect 1392 38596 1448 38598
rect 1680 38106 1736 38108
rect 1760 38106 1816 38108
rect 1680 38054 1690 38106
rect 1690 38054 1736 38106
rect 1760 38054 1806 38106
rect 1806 38054 1816 38106
rect 1680 38052 1736 38054
rect 1760 38052 1816 38054
rect 1312 37562 1368 37564
rect 1392 37562 1448 37564
rect 1312 37510 1322 37562
rect 1322 37510 1368 37562
rect 1392 37510 1438 37562
rect 1438 37510 1448 37562
rect 1312 37508 1368 37510
rect 1392 37508 1448 37510
rect 1680 37018 1736 37020
rect 1760 37018 1816 37020
rect 1680 36966 1690 37018
rect 1690 36966 1736 37018
rect 1760 36966 1806 37018
rect 1806 36966 1816 37018
rect 1680 36964 1736 36966
rect 1760 36964 1816 36966
rect 1312 36474 1368 36476
rect 1392 36474 1448 36476
rect 1312 36422 1322 36474
rect 1322 36422 1368 36474
rect 1392 36422 1438 36474
rect 1438 36422 1448 36474
rect 1312 36420 1368 36422
rect 1392 36420 1448 36422
rect 1680 35930 1736 35932
rect 1760 35930 1816 35932
rect 1680 35878 1690 35930
rect 1690 35878 1736 35930
rect 1760 35878 1806 35930
rect 1806 35878 1816 35930
rect 1680 35876 1736 35878
rect 1760 35876 1816 35878
rect 1312 35386 1368 35388
rect 1392 35386 1448 35388
rect 1312 35334 1322 35386
rect 1322 35334 1368 35386
rect 1392 35334 1438 35386
rect 1438 35334 1448 35386
rect 1312 35332 1368 35334
rect 1392 35332 1448 35334
rect 1680 34842 1736 34844
rect 1760 34842 1816 34844
rect 1680 34790 1690 34842
rect 1690 34790 1736 34842
rect 1760 34790 1806 34842
rect 1806 34790 1816 34842
rect 1680 34788 1736 34790
rect 1760 34788 1816 34790
rect 1312 34298 1368 34300
rect 1392 34298 1448 34300
rect 1312 34246 1322 34298
rect 1322 34246 1368 34298
rect 1392 34246 1438 34298
rect 1438 34246 1448 34298
rect 1312 34244 1368 34246
rect 1392 34244 1448 34246
rect 1680 33754 1736 33756
rect 1760 33754 1816 33756
rect 1680 33702 1690 33754
rect 1690 33702 1736 33754
rect 1760 33702 1806 33754
rect 1806 33702 1816 33754
rect 1680 33700 1736 33702
rect 1760 33700 1816 33702
rect 1312 33210 1368 33212
rect 1392 33210 1448 33212
rect 1312 33158 1322 33210
rect 1322 33158 1368 33210
rect 1392 33158 1438 33210
rect 1438 33158 1448 33210
rect 1312 33156 1368 33158
rect 1392 33156 1448 33158
rect 1680 32666 1736 32668
rect 1760 32666 1816 32668
rect 1680 32614 1690 32666
rect 1690 32614 1736 32666
rect 1760 32614 1806 32666
rect 1806 32614 1816 32666
rect 1680 32612 1736 32614
rect 1760 32612 1816 32614
rect 1312 32122 1368 32124
rect 1392 32122 1448 32124
rect 1312 32070 1322 32122
rect 1322 32070 1368 32122
rect 1392 32070 1438 32122
rect 1438 32070 1448 32122
rect 1312 32068 1368 32070
rect 1392 32068 1448 32070
rect 1680 31578 1736 31580
rect 1760 31578 1816 31580
rect 1680 31526 1690 31578
rect 1690 31526 1736 31578
rect 1760 31526 1806 31578
rect 1806 31526 1816 31578
rect 1680 31524 1736 31526
rect 1760 31524 1816 31526
rect 1312 31034 1368 31036
rect 1392 31034 1448 31036
rect 1312 30982 1322 31034
rect 1322 30982 1368 31034
rect 1392 30982 1438 31034
rect 1438 30982 1448 31034
rect 1312 30980 1368 30982
rect 1392 30980 1448 30982
rect 1680 30490 1736 30492
rect 1760 30490 1816 30492
rect 1680 30438 1690 30490
rect 1690 30438 1736 30490
rect 1760 30438 1806 30490
rect 1806 30438 1816 30490
rect 1680 30436 1736 30438
rect 1760 30436 1816 30438
rect 1312 29946 1368 29948
rect 1392 29946 1448 29948
rect 1312 29894 1322 29946
rect 1322 29894 1368 29946
rect 1392 29894 1438 29946
rect 1438 29894 1448 29946
rect 1312 29892 1368 29894
rect 1392 29892 1448 29894
rect 1680 29402 1736 29404
rect 1760 29402 1816 29404
rect 1680 29350 1690 29402
rect 1690 29350 1736 29402
rect 1760 29350 1806 29402
rect 1806 29350 1816 29402
rect 1680 29348 1736 29350
rect 1760 29348 1816 29350
rect 1312 28858 1368 28860
rect 1392 28858 1448 28860
rect 1312 28806 1322 28858
rect 1322 28806 1368 28858
rect 1392 28806 1438 28858
rect 1438 28806 1448 28858
rect 1312 28804 1368 28806
rect 1392 28804 1448 28806
rect 1680 28314 1736 28316
rect 1760 28314 1816 28316
rect 1680 28262 1690 28314
rect 1690 28262 1736 28314
rect 1760 28262 1806 28314
rect 1806 28262 1816 28314
rect 1680 28260 1736 28262
rect 1760 28260 1816 28262
rect 1312 27770 1368 27772
rect 1392 27770 1448 27772
rect 1312 27718 1322 27770
rect 1322 27718 1368 27770
rect 1392 27718 1438 27770
rect 1438 27718 1448 27770
rect 1312 27716 1368 27718
rect 1392 27716 1448 27718
rect 1680 27226 1736 27228
rect 1760 27226 1816 27228
rect 1680 27174 1690 27226
rect 1690 27174 1736 27226
rect 1760 27174 1806 27226
rect 1806 27174 1816 27226
rect 1680 27172 1736 27174
rect 1760 27172 1816 27174
rect 1312 26682 1368 26684
rect 1392 26682 1448 26684
rect 1312 26630 1322 26682
rect 1322 26630 1368 26682
rect 1392 26630 1438 26682
rect 1438 26630 1448 26682
rect 1312 26628 1368 26630
rect 1392 26628 1448 26630
rect 1680 26138 1736 26140
rect 1760 26138 1816 26140
rect 1680 26086 1690 26138
rect 1690 26086 1736 26138
rect 1760 26086 1806 26138
rect 1806 26086 1816 26138
rect 1680 26084 1736 26086
rect 1760 26084 1816 26086
rect 1312 25594 1368 25596
rect 1392 25594 1448 25596
rect 1312 25542 1322 25594
rect 1322 25542 1368 25594
rect 1392 25542 1438 25594
rect 1438 25542 1448 25594
rect 1312 25540 1368 25542
rect 1392 25540 1448 25542
rect 1680 25050 1736 25052
rect 1760 25050 1816 25052
rect 1680 24998 1690 25050
rect 1690 24998 1736 25050
rect 1760 24998 1806 25050
rect 1806 24998 1816 25050
rect 1680 24996 1736 24998
rect 1760 24996 1816 24998
rect 1312 24506 1368 24508
rect 1392 24506 1448 24508
rect 1312 24454 1322 24506
rect 1322 24454 1368 24506
rect 1392 24454 1438 24506
rect 1438 24454 1448 24506
rect 1312 24452 1368 24454
rect 1392 24452 1448 24454
rect 1680 23962 1736 23964
rect 1760 23962 1816 23964
rect 1680 23910 1690 23962
rect 1690 23910 1736 23962
rect 1760 23910 1806 23962
rect 1806 23910 1816 23962
rect 1680 23908 1736 23910
rect 1760 23908 1816 23910
rect 1312 23418 1368 23420
rect 1392 23418 1448 23420
rect 1312 23366 1322 23418
rect 1322 23366 1368 23418
rect 1392 23366 1438 23418
rect 1438 23366 1448 23418
rect 1312 23364 1368 23366
rect 1392 23364 1448 23366
rect 1680 22874 1736 22876
rect 1760 22874 1816 22876
rect 1680 22822 1690 22874
rect 1690 22822 1736 22874
rect 1760 22822 1806 22874
rect 1806 22822 1816 22874
rect 1680 22820 1736 22822
rect 1760 22820 1816 22822
rect 1312 22330 1368 22332
rect 1392 22330 1448 22332
rect 1312 22278 1322 22330
rect 1322 22278 1368 22330
rect 1392 22278 1438 22330
rect 1438 22278 1448 22330
rect 1312 22276 1368 22278
rect 1392 22276 1448 22278
rect 1680 21786 1736 21788
rect 1760 21786 1816 21788
rect 1680 21734 1690 21786
rect 1690 21734 1736 21786
rect 1760 21734 1806 21786
rect 1806 21734 1816 21786
rect 1680 21732 1736 21734
rect 1760 21732 1816 21734
rect 1312 21242 1368 21244
rect 1392 21242 1448 21244
rect 1312 21190 1322 21242
rect 1322 21190 1368 21242
rect 1392 21190 1438 21242
rect 1438 21190 1448 21242
rect 1312 21188 1368 21190
rect 1392 21188 1448 21190
rect 1680 20698 1736 20700
rect 1760 20698 1816 20700
rect 1680 20646 1690 20698
rect 1690 20646 1736 20698
rect 1760 20646 1806 20698
rect 1806 20646 1816 20698
rect 1680 20644 1736 20646
rect 1760 20644 1816 20646
rect 1312 20154 1368 20156
rect 1392 20154 1448 20156
rect 1312 20102 1322 20154
rect 1322 20102 1368 20154
rect 1392 20102 1438 20154
rect 1438 20102 1448 20154
rect 1312 20100 1368 20102
rect 1392 20100 1448 20102
rect 1680 19610 1736 19612
rect 1760 19610 1816 19612
rect 1680 19558 1690 19610
rect 1690 19558 1736 19610
rect 1760 19558 1806 19610
rect 1806 19558 1816 19610
rect 1680 19556 1736 19558
rect 1760 19556 1816 19558
rect 1312 19066 1368 19068
rect 1392 19066 1448 19068
rect 1312 19014 1322 19066
rect 1322 19014 1368 19066
rect 1392 19014 1438 19066
rect 1438 19014 1448 19066
rect 1312 19012 1368 19014
rect 1392 19012 1448 19014
rect 1680 18522 1736 18524
rect 1760 18522 1816 18524
rect 1680 18470 1690 18522
rect 1690 18470 1736 18522
rect 1760 18470 1806 18522
rect 1806 18470 1816 18522
rect 1680 18468 1736 18470
rect 1760 18468 1816 18470
rect 1312 17978 1368 17980
rect 1392 17978 1448 17980
rect 1312 17926 1322 17978
rect 1322 17926 1368 17978
rect 1392 17926 1438 17978
rect 1438 17926 1448 17978
rect 1312 17924 1368 17926
rect 1392 17924 1448 17926
rect 1680 17434 1736 17436
rect 1760 17434 1816 17436
rect 1680 17382 1690 17434
rect 1690 17382 1736 17434
rect 1760 17382 1806 17434
rect 1806 17382 1816 17434
rect 1680 17380 1736 17382
rect 1760 17380 1816 17382
rect 1312 16890 1368 16892
rect 1392 16890 1448 16892
rect 1312 16838 1322 16890
rect 1322 16838 1368 16890
rect 1392 16838 1438 16890
rect 1438 16838 1448 16890
rect 1312 16836 1368 16838
rect 1392 16836 1448 16838
rect 1680 16346 1736 16348
rect 1760 16346 1816 16348
rect 1680 16294 1690 16346
rect 1690 16294 1736 16346
rect 1760 16294 1806 16346
rect 1806 16294 1816 16346
rect 1680 16292 1736 16294
rect 1760 16292 1816 16294
rect 1312 15802 1368 15804
rect 1392 15802 1448 15804
rect 1312 15750 1322 15802
rect 1322 15750 1368 15802
rect 1392 15750 1438 15802
rect 1438 15750 1448 15802
rect 1312 15748 1368 15750
rect 1392 15748 1448 15750
rect 1680 15258 1736 15260
rect 1760 15258 1816 15260
rect 1680 15206 1690 15258
rect 1690 15206 1736 15258
rect 1760 15206 1806 15258
rect 1806 15206 1816 15258
rect 1680 15204 1736 15206
rect 1760 15204 1816 15206
rect 1312 14714 1368 14716
rect 1392 14714 1448 14716
rect 1312 14662 1322 14714
rect 1322 14662 1368 14714
rect 1392 14662 1438 14714
rect 1438 14662 1448 14714
rect 1312 14660 1368 14662
rect 1392 14660 1448 14662
rect 1680 14170 1736 14172
rect 1760 14170 1816 14172
rect 1680 14118 1690 14170
rect 1690 14118 1736 14170
rect 1760 14118 1806 14170
rect 1806 14118 1816 14170
rect 1680 14116 1736 14118
rect 1760 14116 1816 14118
rect 1312 13626 1368 13628
rect 1392 13626 1448 13628
rect 1312 13574 1322 13626
rect 1322 13574 1368 13626
rect 1392 13574 1438 13626
rect 1438 13574 1448 13626
rect 1312 13572 1368 13574
rect 1392 13572 1448 13574
rect 1680 13082 1736 13084
rect 1760 13082 1816 13084
rect 1680 13030 1690 13082
rect 1690 13030 1736 13082
rect 1760 13030 1806 13082
rect 1806 13030 1816 13082
rect 1680 13028 1736 13030
rect 1760 13028 1816 13030
rect 1312 12538 1368 12540
rect 1392 12538 1448 12540
rect 1312 12486 1322 12538
rect 1322 12486 1368 12538
rect 1392 12486 1438 12538
rect 1438 12486 1448 12538
rect 1312 12484 1368 12486
rect 1392 12484 1448 12486
rect 1680 11994 1736 11996
rect 1760 11994 1816 11996
rect 1680 11942 1690 11994
rect 1690 11942 1736 11994
rect 1760 11942 1806 11994
rect 1806 11942 1816 11994
rect 1680 11940 1736 11942
rect 1760 11940 1816 11942
rect 1312 11450 1368 11452
rect 1392 11450 1448 11452
rect 1312 11398 1322 11450
rect 1322 11398 1368 11450
rect 1392 11398 1438 11450
rect 1438 11398 1448 11450
rect 1312 11396 1368 11398
rect 1392 11396 1448 11398
rect 1680 10906 1736 10908
rect 1760 10906 1816 10908
rect 1680 10854 1690 10906
rect 1690 10854 1736 10906
rect 1760 10854 1806 10906
rect 1806 10854 1816 10906
rect 1680 10852 1736 10854
rect 1760 10852 1816 10854
rect 1312 10362 1368 10364
rect 1392 10362 1448 10364
rect 1312 10310 1322 10362
rect 1322 10310 1368 10362
rect 1392 10310 1438 10362
rect 1438 10310 1448 10362
rect 1312 10308 1368 10310
rect 1392 10308 1448 10310
rect 1680 9818 1736 9820
rect 1760 9818 1816 9820
rect 1680 9766 1690 9818
rect 1690 9766 1736 9818
rect 1760 9766 1806 9818
rect 1806 9766 1816 9818
rect 1680 9764 1736 9766
rect 1760 9764 1816 9766
rect 1312 9274 1368 9276
rect 1392 9274 1448 9276
rect 1312 9222 1322 9274
rect 1322 9222 1368 9274
rect 1392 9222 1438 9274
rect 1438 9222 1448 9274
rect 1312 9220 1368 9222
rect 1392 9220 1448 9222
rect 1680 8730 1736 8732
rect 1760 8730 1816 8732
rect 1680 8678 1690 8730
rect 1690 8678 1736 8730
rect 1760 8678 1806 8730
rect 1806 8678 1816 8730
rect 1680 8676 1736 8678
rect 1760 8676 1816 8678
rect 1312 8186 1368 8188
rect 1392 8186 1448 8188
rect 1312 8134 1322 8186
rect 1322 8134 1368 8186
rect 1392 8134 1438 8186
rect 1438 8134 1448 8186
rect 1312 8132 1368 8134
rect 1392 8132 1448 8134
rect 1680 7642 1736 7644
rect 1760 7642 1816 7644
rect 1680 7590 1690 7642
rect 1690 7590 1736 7642
rect 1760 7590 1806 7642
rect 1806 7590 1816 7642
rect 1680 7588 1736 7590
rect 1760 7588 1816 7590
rect 1312 7098 1368 7100
rect 1392 7098 1448 7100
rect 1312 7046 1322 7098
rect 1322 7046 1368 7098
rect 1392 7046 1438 7098
rect 1438 7046 1448 7098
rect 1312 7044 1368 7046
rect 1392 7044 1448 7046
rect 1680 6554 1736 6556
rect 1760 6554 1816 6556
rect 1680 6502 1690 6554
rect 1690 6502 1736 6554
rect 1760 6502 1806 6554
rect 1806 6502 1816 6554
rect 1680 6500 1736 6502
rect 1760 6500 1816 6502
rect 1312 6010 1368 6012
rect 1392 6010 1448 6012
rect 1312 5958 1322 6010
rect 1322 5958 1368 6010
rect 1392 5958 1438 6010
rect 1438 5958 1448 6010
rect 1312 5956 1368 5958
rect 1392 5956 1448 5958
rect 1680 5466 1736 5468
rect 1760 5466 1816 5468
rect 1680 5414 1690 5466
rect 1690 5414 1736 5466
rect 1760 5414 1806 5466
rect 1806 5414 1816 5466
rect 1680 5412 1736 5414
rect 1760 5412 1816 5414
rect 1312 4922 1368 4924
rect 1392 4922 1448 4924
rect 1312 4870 1322 4922
rect 1322 4870 1368 4922
rect 1392 4870 1438 4922
rect 1438 4870 1448 4922
rect 1312 4868 1368 4870
rect 1392 4868 1448 4870
rect 1680 4378 1736 4380
rect 1760 4378 1816 4380
rect 1680 4326 1690 4378
rect 1690 4326 1736 4378
rect 1760 4326 1806 4378
rect 1806 4326 1816 4378
rect 1680 4324 1736 4326
rect 1760 4324 1816 4326
rect 35600 60954 35656 60956
rect 35680 60954 35736 60956
rect 35760 60954 35816 60956
rect 35840 60954 35896 60956
rect 35600 60902 35646 60954
rect 35646 60902 35656 60954
rect 35680 60902 35710 60954
rect 35710 60902 35722 60954
rect 35722 60902 35736 60954
rect 35760 60902 35774 60954
rect 35774 60902 35786 60954
rect 35786 60902 35816 60954
rect 35840 60902 35850 60954
rect 35850 60902 35896 60954
rect 35600 60900 35656 60902
rect 35680 60900 35736 60902
rect 35760 60900 35816 60902
rect 35840 60900 35896 60902
rect 66320 101210 66376 101212
rect 66400 101210 66456 101212
rect 66480 101210 66536 101212
rect 66560 101210 66616 101212
rect 66320 101158 66366 101210
rect 66366 101158 66376 101210
rect 66400 101158 66430 101210
rect 66430 101158 66442 101210
rect 66442 101158 66456 101210
rect 66480 101158 66494 101210
rect 66494 101158 66506 101210
rect 66506 101158 66536 101210
rect 66560 101158 66570 101210
rect 66570 101158 66616 101210
rect 66320 101156 66376 101158
rect 66400 101156 66456 101158
rect 66480 101156 66536 101158
rect 66560 101156 66616 101158
rect 97040 101210 97096 101212
rect 97120 101210 97176 101212
rect 97200 101210 97256 101212
rect 97280 101210 97336 101212
rect 97040 101158 97086 101210
rect 97086 101158 97096 101210
rect 97120 101158 97150 101210
rect 97150 101158 97162 101210
rect 97162 101158 97176 101210
rect 97200 101158 97214 101210
rect 97214 101158 97226 101210
rect 97226 101158 97256 101210
rect 97280 101158 97290 101210
rect 97290 101158 97336 101210
rect 97040 101156 97096 101158
rect 97120 101156 97176 101158
rect 97200 101156 97256 101158
rect 97280 101156 97336 101158
rect 65660 100666 65716 100668
rect 65740 100666 65796 100668
rect 65820 100666 65876 100668
rect 65900 100666 65956 100668
rect 65660 100614 65706 100666
rect 65706 100614 65716 100666
rect 65740 100614 65770 100666
rect 65770 100614 65782 100666
rect 65782 100614 65796 100666
rect 65820 100614 65834 100666
rect 65834 100614 65846 100666
rect 65846 100614 65876 100666
rect 65900 100614 65910 100666
rect 65910 100614 65956 100666
rect 65660 100612 65716 100614
rect 65740 100612 65796 100614
rect 65820 100612 65876 100614
rect 65900 100612 65956 100614
rect 96380 100666 96436 100668
rect 96460 100666 96516 100668
rect 96540 100666 96596 100668
rect 96620 100666 96676 100668
rect 96380 100614 96426 100666
rect 96426 100614 96436 100666
rect 96460 100614 96490 100666
rect 96490 100614 96502 100666
rect 96502 100614 96516 100666
rect 96540 100614 96554 100666
rect 96554 100614 96566 100666
rect 96566 100614 96596 100666
rect 96620 100614 96630 100666
rect 96630 100614 96676 100666
rect 96380 100612 96436 100614
rect 96460 100612 96516 100614
rect 96540 100612 96596 100614
rect 96620 100612 96676 100614
rect 66320 100122 66376 100124
rect 66400 100122 66456 100124
rect 66480 100122 66536 100124
rect 66560 100122 66616 100124
rect 66320 100070 66366 100122
rect 66366 100070 66376 100122
rect 66400 100070 66430 100122
rect 66430 100070 66442 100122
rect 66442 100070 66456 100122
rect 66480 100070 66494 100122
rect 66494 100070 66506 100122
rect 66506 100070 66536 100122
rect 66560 100070 66570 100122
rect 66570 100070 66616 100122
rect 66320 100068 66376 100070
rect 66400 100068 66456 100070
rect 66480 100068 66536 100070
rect 66560 100068 66616 100070
rect 97040 100122 97096 100124
rect 97120 100122 97176 100124
rect 97200 100122 97256 100124
rect 97280 100122 97336 100124
rect 97040 100070 97086 100122
rect 97086 100070 97096 100122
rect 97120 100070 97150 100122
rect 97150 100070 97162 100122
rect 97162 100070 97176 100122
rect 97200 100070 97214 100122
rect 97214 100070 97226 100122
rect 97226 100070 97256 100122
rect 97280 100070 97290 100122
rect 97290 100070 97336 100122
rect 97040 100068 97096 100070
rect 97120 100068 97176 100070
rect 97200 100068 97256 100070
rect 97280 100068 97336 100070
rect 65660 99578 65716 99580
rect 65740 99578 65796 99580
rect 65820 99578 65876 99580
rect 65900 99578 65956 99580
rect 65660 99526 65706 99578
rect 65706 99526 65716 99578
rect 65740 99526 65770 99578
rect 65770 99526 65782 99578
rect 65782 99526 65796 99578
rect 65820 99526 65834 99578
rect 65834 99526 65846 99578
rect 65846 99526 65876 99578
rect 65900 99526 65910 99578
rect 65910 99526 65956 99578
rect 65660 99524 65716 99526
rect 65740 99524 65796 99526
rect 65820 99524 65876 99526
rect 65900 99524 65956 99526
rect 96380 99578 96436 99580
rect 96460 99578 96516 99580
rect 96540 99578 96596 99580
rect 96620 99578 96676 99580
rect 96380 99526 96426 99578
rect 96426 99526 96436 99578
rect 96460 99526 96490 99578
rect 96490 99526 96502 99578
rect 96502 99526 96516 99578
rect 96540 99526 96554 99578
rect 96554 99526 96566 99578
rect 96566 99526 96596 99578
rect 96620 99526 96630 99578
rect 96630 99526 96676 99578
rect 96380 99524 96436 99526
rect 96460 99524 96516 99526
rect 96540 99524 96596 99526
rect 96620 99524 96676 99526
rect 66320 99034 66376 99036
rect 66400 99034 66456 99036
rect 66480 99034 66536 99036
rect 66560 99034 66616 99036
rect 66320 98982 66366 99034
rect 66366 98982 66376 99034
rect 66400 98982 66430 99034
rect 66430 98982 66442 99034
rect 66442 98982 66456 99034
rect 66480 98982 66494 99034
rect 66494 98982 66506 99034
rect 66506 98982 66536 99034
rect 66560 98982 66570 99034
rect 66570 98982 66616 99034
rect 66320 98980 66376 98982
rect 66400 98980 66456 98982
rect 66480 98980 66536 98982
rect 66560 98980 66616 98982
rect 97040 99034 97096 99036
rect 97120 99034 97176 99036
rect 97200 99034 97256 99036
rect 97280 99034 97336 99036
rect 97040 98982 97086 99034
rect 97086 98982 97096 99034
rect 97120 98982 97150 99034
rect 97150 98982 97162 99034
rect 97162 98982 97176 99034
rect 97200 98982 97214 99034
rect 97214 98982 97226 99034
rect 97226 98982 97256 99034
rect 97280 98982 97290 99034
rect 97290 98982 97336 99034
rect 97040 98980 97096 98982
rect 97120 98980 97176 98982
rect 97200 98980 97256 98982
rect 97280 98980 97336 98982
rect 65660 98490 65716 98492
rect 65740 98490 65796 98492
rect 65820 98490 65876 98492
rect 65900 98490 65956 98492
rect 65660 98438 65706 98490
rect 65706 98438 65716 98490
rect 65740 98438 65770 98490
rect 65770 98438 65782 98490
rect 65782 98438 65796 98490
rect 65820 98438 65834 98490
rect 65834 98438 65846 98490
rect 65846 98438 65876 98490
rect 65900 98438 65910 98490
rect 65910 98438 65956 98490
rect 65660 98436 65716 98438
rect 65740 98436 65796 98438
rect 65820 98436 65876 98438
rect 65900 98436 65956 98438
rect 96380 98490 96436 98492
rect 96460 98490 96516 98492
rect 96540 98490 96596 98492
rect 96620 98490 96676 98492
rect 96380 98438 96426 98490
rect 96426 98438 96436 98490
rect 96460 98438 96490 98490
rect 96490 98438 96502 98490
rect 96502 98438 96516 98490
rect 96540 98438 96554 98490
rect 96554 98438 96566 98490
rect 96566 98438 96596 98490
rect 96620 98438 96630 98490
rect 96630 98438 96676 98490
rect 96380 98436 96436 98438
rect 96460 98436 96516 98438
rect 96540 98436 96596 98438
rect 96620 98436 96676 98438
rect 66320 97946 66376 97948
rect 66400 97946 66456 97948
rect 66480 97946 66536 97948
rect 66560 97946 66616 97948
rect 66320 97894 66366 97946
rect 66366 97894 66376 97946
rect 66400 97894 66430 97946
rect 66430 97894 66442 97946
rect 66442 97894 66456 97946
rect 66480 97894 66494 97946
rect 66494 97894 66506 97946
rect 66506 97894 66536 97946
rect 66560 97894 66570 97946
rect 66570 97894 66616 97946
rect 66320 97892 66376 97894
rect 66400 97892 66456 97894
rect 66480 97892 66536 97894
rect 66560 97892 66616 97894
rect 97040 97946 97096 97948
rect 97120 97946 97176 97948
rect 97200 97946 97256 97948
rect 97280 97946 97336 97948
rect 97040 97894 97086 97946
rect 97086 97894 97096 97946
rect 97120 97894 97150 97946
rect 97150 97894 97162 97946
rect 97162 97894 97176 97946
rect 97200 97894 97214 97946
rect 97214 97894 97226 97946
rect 97226 97894 97256 97946
rect 97280 97894 97290 97946
rect 97290 97894 97336 97946
rect 97040 97892 97096 97894
rect 97120 97892 97176 97894
rect 97200 97892 97256 97894
rect 97280 97892 97336 97894
rect 65660 97402 65716 97404
rect 65740 97402 65796 97404
rect 65820 97402 65876 97404
rect 65900 97402 65956 97404
rect 65660 97350 65706 97402
rect 65706 97350 65716 97402
rect 65740 97350 65770 97402
rect 65770 97350 65782 97402
rect 65782 97350 65796 97402
rect 65820 97350 65834 97402
rect 65834 97350 65846 97402
rect 65846 97350 65876 97402
rect 65900 97350 65910 97402
rect 65910 97350 65956 97402
rect 65660 97348 65716 97350
rect 65740 97348 65796 97350
rect 65820 97348 65876 97350
rect 65900 97348 65956 97350
rect 96380 97402 96436 97404
rect 96460 97402 96516 97404
rect 96540 97402 96596 97404
rect 96620 97402 96676 97404
rect 96380 97350 96426 97402
rect 96426 97350 96436 97402
rect 96460 97350 96490 97402
rect 96490 97350 96502 97402
rect 96502 97350 96516 97402
rect 96540 97350 96554 97402
rect 96554 97350 96566 97402
rect 96566 97350 96596 97402
rect 96620 97350 96630 97402
rect 96630 97350 96676 97402
rect 96380 97348 96436 97350
rect 96460 97348 96516 97350
rect 96540 97348 96596 97350
rect 96620 97348 96676 97350
rect 66320 96858 66376 96860
rect 66400 96858 66456 96860
rect 66480 96858 66536 96860
rect 66560 96858 66616 96860
rect 66320 96806 66366 96858
rect 66366 96806 66376 96858
rect 66400 96806 66430 96858
rect 66430 96806 66442 96858
rect 66442 96806 66456 96858
rect 66480 96806 66494 96858
rect 66494 96806 66506 96858
rect 66506 96806 66536 96858
rect 66560 96806 66570 96858
rect 66570 96806 66616 96858
rect 66320 96804 66376 96806
rect 66400 96804 66456 96806
rect 66480 96804 66536 96806
rect 66560 96804 66616 96806
rect 97040 96858 97096 96860
rect 97120 96858 97176 96860
rect 97200 96858 97256 96860
rect 97280 96858 97336 96860
rect 97040 96806 97086 96858
rect 97086 96806 97096 96858
rect 97120 96806 97150 96858
rect 97150 96806 97162 96858
rect 97162 96806 97176 96858
rect 97200 96806 97214 96858
rect 97214 96806 97226 96858
rect 97226 96806 97256 96858
rect 97280 96806 97290 96858
rect 97290 96806 97336 96858
rect 97040 96804 97096 96806
rect 97120 96804 97176 96806
rect 97200 96804 97256 96806
rect 97280 96804 97336 96806
rect 65660 96314 65716 96316
rect 65740 96314 65796 96316
rect 65820 96314 65876 96316
rect 65900 96314 65956 96316
rect 65660 96262 65706 96314
rect 65706 96262 65716 96314
rect 65740 96262 65770 96314
rect 65770 96262 65782 96314
rect 65782 96262 65796 96314
rect 65820 96262 65834 96314
rect 65834 96262 65846 96314
rect 65846 96262 65876 96314
rect 65900 96262 65910 96314
rect 65910 96262 65956 96314
rect 65660 96260 65716 96262
rect 65740 96260 65796 96262
rect 65820 96260 65876 96262
rect 65900 96260 65956 96262
rect 96380 96314 96436 96316
rect 96460 96314 96516 96316
rect 96540 96314 96596 96316
rect 96620 96314 96676 96316
rect 96380 96262 96426 96314
rect 96426 96262 96436 96314
rect 96460 96262 96490 96314
rect 96490 96262 96502 96314
rect 96502 96262 96516 96314
rect 96540 96262 96554 96314
rect 96554 96262 96566 96314
rect 96566 96262 96596 96314
rect 96620 96262 96630 96314
rect 96630 96262 96676 96314
rect 96380 96260 96436 96262
rect 96460 96260 96516 96262
rect 96540 96260 96596 96262
rect 96620 96260 96676 96262
rect 66320 95770 66376 95772
rect 66400 95770 66456 95772
rect 66480 95770 66536 95772
rect 66560 95770 66616 95772
rect 66320 95718 66366 95770
rect 66366 95718 66376 95770
rect 66400 95718 66430 95770
rect 66430 95718 66442 95770
rect 66442 95718 66456 95770
rect 66480 95718 66494 95770
rect 66494 95718 66506 95770
rect 66506 95718 66536 95770
rect 66560 95718 66570 95770
rect 66570 95718 66616 95770
rect 66320 95716 66376 95718
rect 66400 95716 66456 95718
rect 66480 95716 66536 95718
rect 66560 95716 66616 95718
rect 97040 95770 97096 95772
rect 97120 95770 97176 95772
rect 97200 95770 97256 95772
rect 97280 95770 97336 95772
rect 97040 95718 97086 95770
rect 97086 95718 97096 95770
rect 97120 95718 97150 95770
rect 97150 95718 97162 95770
rect 97162 95718 97176 95770
rect 97200 95718 97214 95770
rect 97214 95718 97226 95770
rect 97226 95718 97256 95770
rect 97280 95718 97290 95770
rect 97290 95718 97336 95770
rect 97040 95716 97096 95718
rect 97120 95716 97176 95718
rect 97200 95716 97256 95718
rect 97280 95716 97336 95718
rect 65660 95226 65716 95228
rect 65740 95226 65796 95228
rect 65820 95226 65876 95228
rect 65900 95226 65956 95228
rect 65660 95174 65706 95226
rect 65706 95174 65716 95226
rect 65740 95174 65770 95226
rect 65770 95174 65782 95226
rect 65782 95174 65796 95226
rect 65820 95174 65834 95226
rect 65834 95174 65846 95226
rect 65846 95174 65876 95226
rect 65900 95174 65910 95226
rect 65910 95174 65956 95226
rect 65660 95172 65716 95174
rect 65740 95172 65796 95174
rect 65820 95172 65876 95174
rect 65900 95172 65956 95174
rect 96380 95226 96436 95228
rect 96460 95226 96516 95228
rect 96540 95226 96596 95228
rect 96620 95226 96676 95228
rect 96380 95174 96426 95226
rect 96426 95174 96436 95226
rect 96460 95174 96490 95226
rect 96490 95174 96502 95226
rect 96502 95174 96516 95226
rect 96540 95174 96554 95226
rect 96554 95174 96566 95226
rect 96566 95174 96596 95226
rect 96620 95174 96630 95226
rect 96630 95174 96676 95226
rect 96380 95172 96436 95174
rect 96460 95172 96516 95174
rect 96540 95172 96596 95174
rect 96620 95172 96676 95174
rect 66320 94682 66376 94684
rect 66400 94682 66456 94684
rect 66480 94682 66536 94684
rect 66560 94682 66616 94684
rect 66320 94630 66366 94682
rect 66366 94630 66376 94682
rect 66400 94630 66430 94682
rect 66430 94630 66442 94682
rect 66442 94630 66456 94682
rect 66480 94630 66494 94682
rect 66494 94630 66506 94682
rect 66506 94630 66536 94682
rect 66560 94630 66570 94682
rect 66570 94630 66616 94682
rect 66320 94628 66376 94630
rect 66400 94628 66456 94630
rect 66480 94628 66536 94630
rect 66560 94628 66616 94630
rect 97040 94682 97096 94684
rect 97120 94682 97176 94684
rect 97200 94682 97256 94684
rect 97280 94682 97336 94684
rect 97040 94630 97086 94682
rect 97086 94630 97096 94682
rect 97120 94630 97150 94682
rect 97150 94630 97162 94682
rect 97162 94630 97176 94682
rect 97200 94630 97214 94682
rect 97214 94630 97226 94682
rect 97226 94630 97256 94682
rect 97280 94630 97290 94682
rect 97290 94630 97336 94682
rect 97040 94628 97096 94630
rect 97120 94628 97176 94630
rect 97200 94628 97256 94630
rect 97280 94628 97336 94630
rect 65660 94138 65716 94140
rect 65740 94138 65796 94140
rect 65820 94138 65876 94140
rect 65900 94138 65956 94140
rect 65660 94086 65706 94138
rect 65706 94086 65716 94138
rect 65740 94086 65770 94138
rect 65770 94086 65782 94138
rect 65782 94086 65796 94138
rect 65820 94086 65834 94138
rect 65834 94086 65846 94138
rect 65846 94086 65876 94138
rect 65900 94086 65910 94138
rect 65910 94086 65956 94138
rect 65660 94084 65716 94086
rect 65740 94084 65796 94086
rect 65820 94084 65876 94086
rect 65900 94084 65956 94086
rect 96380 94138 96436 94140
rect 96460 94138 96516 94140
rect 96540 94138 96596 94140
rect 96620 94138 96676 94140
rect 96380 94086 96426 94138
rect 96426 94086 96436 94138
rect 96460 94086 96490 94138
rect 96490 94086 96502 94138
rect 96502 94086 96516 94138
rect 96540 94086 96554 94138
rect 96554 94086 96566 94138
rect 96566 94086 96596 94138
rect 96620 94086 96630 94138
rect 96630 94086 96676 94138
rect 96380 94084 96436 94086
rect 96460 94084 96516 94086
rect 96540 94084 96596 94086
rect 96620 94084 96676 94086
rect 66320 93594 66376 93596
rect 66400 93594 66456 93596
rect 66480 93594 66536 93596
rect 66560 93594 66616 93596
rect 66320 93542 66366 93594
rect 66366 93542 66376 93594
rect 66400 93542 66430 93594
rect 66430 93542 66442 93594
rect 66442 93542 66456 93594
rect 66480 93542 66494 93594
rect 66494 93542 66506 93594
rect 66506 93542 66536 93594
rect 66560 93542 66570 93594
rect 66570 93542 66616 93594
rect 66320 93540 66376 93542
rect 66400 93540 66456 93542
rect 66480 93540 66536 93542
rect 66560 93540 66616 93542
rect 97040 93594 97096 93596
rect 97120 93594 97176 93596
rect 97200 93594 97256 93596
rect 97280 93594 97336 93596
rect 97040 93542 97086 93594
rect 97086 93542 97096 93594
rect 97120 93542 97150 93594
rect 97150 93542 97162 93594
rect 97162 93542 97176 93594
rect 97200 93542 97214 93594
rect 97214 93542 97226 93594
rect 97226 93542 97256 93594
rect 97280 93542 97290 93594
rect 97290 93542 97336 93594
rect 97040 93540 97096 93542
rect 97120 93540 97176 93542
rect 97200 93540 97256 93542
rect 97280 93540 97336 93542
rect 65660 93050 65716 93052
rect 65740 93050 65796 93052
rect 65820 93050 65876 93052
rect 65900 93050 65956 93052
rect 65660 92998 65706 93050
rect 65706 92998 65716 93050
rect 65740 92998 65770 93050
rect 65770 92998 65782 93050
rect 65782 92998 65796 93050
rect 65820 92998 65834 93050
rect 65834 92998 65846 93050
rect 65846 92998 65876 93050
rect 65900 92998 65910 93050
rect 65910 92998 65956 93050
rect 65660 92996 65716 92998
rect 65740 92996 65796 92998
rect 65820 92996 65876 92998
rect 65900 92996 65956 92998
rect 96380 93050 96436 93052
rect 96460 93050 96516 93052
rect 96540 93050 96596 93052
rect 96620 93050 96676 93052
rect 96380 92998 96426 93050
rect 96426 92998 96436 93050
rect 96460 92998 96490 93050
rect 96490 92998 96502 93050
rect 96502 92998 96516 93050
rect 96540 92998 96554 93050
rect 96554 92998 96566 93050
rect 96566 92998 96596 93050
rect 96620 92998 96630 93050
rect 96630 92998 96676 93050
rect 96380 92996 96436 92998
rect 96460 92996 96516 92998
rect 96540 92996 96596 92998
rect 96620 92996 96676 92998
rect 66320 92506 66376 92508
rect 66400 92506 66456 92508
rect 66480 92506 66536 92508
rect 66560 92506 66616 92508
rect 66320 92454 66366 92506
rect 66366 92454 66376 92506
rect 66400 92454 66430 92506
rect 66430 92454 66442 92506
rect 66442 92454 66456 92506
rect 66480 92454 66494 92506
rect 66494 92454 66506 92506
rect 66506 92454 66536 92506
rect 66560 92454 66570 92506
rect 66570 92454 66616 92506
rect 66320 92452 66376 92454
rect 66400 92452 66456 92454
rect 66480 92452 66536 92454
rect 66560 92452 66616 92454
rect 97040 92506 97096 92508
rect 97120 92506 97176 92508
rect 97200 92506 97256 92508
rect 97280 92506 97336 92508
rect 97040 92454 97086 92506
rect 97086 92454 97096 92506
rect 97120 92454 97150 92506
rect 97150 92454 97162 92506
rect 97162 92454 97176 92506
rect 97200 92454 97214 92506
rect 97214 92454 97226 92506
rect 97226 92454 97256 92506
rect 97280 92454 97290 92506
rect 97290 92454 97336 92506
rect 97040 92452 97096 92454
rect 97120 92452 97176 92454
rect 97200 92452 97256 92454
rect 97280 92452 97336 92454
rect 65660 91962 65716 91964
rect 65740 91962 65796 91964
rect 65820 91962 65876 91964
rect 65900 91962 65956 91964
rect 65660 91910 65706 91962
rect 65706 91910 65716 91962
rect 65740 91910 65770 91962
rect 65770 91910 65782 91962
rect 65782 91910 65796 91962
rect 65820 91910 65834 91962
rect 65834 91910 65846 91962
rect 65846 91910 65876 91962
rect 65900 91910 65910 91962
rect 65910 91910 65956 91962
rect 65660 91908 65716 91910
rect 65740 91908 65796 91910
rect 65820 91908 65876 91910
rect 65900 91908 65956 91910
rect 96380 91962 96436 91964
rect 96460 91962 96516 91964
rect 96540 91962 96596 91964
rect 96620 91962 96676 91964
rect 96380 91910 96426 91962
rect 96426 91910 96436 91962
rect 96460 91910 96490 91962
rect 96490 91910 96502 91962
rect 96502 91910 96516 91962
rect 96540 91910 96554 91962
rect 96554 91910 96566 91962
rect 96566 91910 96596 91962
rect 96620 91910 96630 91962
rect 96630 91910 96676 91962
rect 96380 91908 96436 91910
rect 96460 91908 96516 91910
rect 96540 91908 96596 91910
rect 96620 91908 96676 91910
rect 66320 91418 66376 91420
rect 66400 91418 66456 91420
rect 66480 91418 66536 91420
rect 66560 91418 66616 91420
rect 66320 91366 66366 91418
rect 66366 91366 66376 91418
rect 66400 91366 66430 91418
rect 66430 91366 66442 91418
rect 66442 91366 66456 91418
rect 66480 91366 66494 91418
rect 66494 91366 66506 91418
rect 66506 91366 66536 91418
rect 66560 91366 66570 91418
rect 66570 91366 66616 91418
rect 66320 91364 66376 91366
rect 66400 91364 66456 91366
rect 66480 91364 66536 91366
rect 66560 91364 66616 91366
rect 97040 91418 97096 91420
rect 97120 91418 97176 91420
rect 97200 91418 97256 91420
rect 97280 91418 97336 91420
rect 97040 91366 97086 91418
rect 97086 91366 97096 91418
rect 97120 91366 97150 91418
rect 97150 91366 97162 91418
rect 97162 91366 97176 91418
rect 97200 91366 97214 91418
rect 97214 91366 97226 91418
rect 97226 91366 97256 91418
rect 97280 91366 97290 91418
rect 97290 91366 97336 91418
rect 97040 91364 97096 91366
rect 97120 91364 97176 91366
rect 97200 91364 97256 91366
rect 97280 91364 97336 91366
rect 65660 90874 65716 90876
rect 65740 90874 65796 90876
rect 65820 90874 65876 90876
rect 65900 90874 65956 90876
rect 65660 90822 65706 90874
rect 65706 90822 65716 90874
rect 65740 90822 65770 90874
rect 65770 90822 65782 90874
rect 65782 90822 65796 90874
rect 65820 90822 65834 90874
rect 65834 90822 65846 90874
rect 65846 90822 65876 90874
rect 65900 90822 65910 90874
rect 65910 90822 65956 90874
rect 65660 90820 65716 90822
rect 65740 90820 65796 90822
rect 65820 90820 65876 90822
rect 65900 90820 65956 90822
rect 96380 90874 96436 90876
rect 96460 90874 96516 90876
rect 96540 90874 96596 90876
rect 96620 90874 96676 90876
rect 96380 90822 96426 90874
rect 96426 90822 96436 90874
rect 96460 90822 96490 90874
rect 96490 90822 96502 90874
rect 96502 90822 96516 90874
rect 96540 90822 96554 90874
rect 96554 90822 96566 90874
rect 96566 90822 96596 90874
rect 96620 90822 96630 90874
rect 96630 90822 96676 90874
rect 96380 90820 96436 90822
rect 96460 90820 96516 90822
rect 96540 90820 96596 90822
rect 96620 90820 96676 90822
rect 66320 90330 66376 90332
rect 66400 90330 66456 90332
rect 66480 90330 66536 90332
rect 66560 90330 66616 90332
rect 66320 90278 66366 90330
rect 66366 90278 66376 90330
rect 66400 90278 66430 90330
rect 66430 90278 66442 90330
rect 66442 90278 66456 90330
rect 66480 90278 66494 90330
rect 66494 90278 66506 90330
rect 66506 90278 66536 90330
rect 66560 90278 66570 90330
rect 66570 90278 66616 90330
rect 66320 90276 66376 90278
rect 66400 90276 66456 90278
rect 66480 90276 66536 90278
rect 66560 90276 66616 90278
rect 97040 90330 97096 90332
rect 97120 90330 97176 90332
rect 97200 90330 97256 90332
rect 97280 90330 97336 90332
rect 97040 90278 97086 90330
rect 97086 90278 97096 90330
rect 97120 90278 97150 90330
rect 97150 90278 97162 90330
rect 97162 90278 97176 90330
rect 97200 90278 97214 90330
rect 97214 90278 97226 90330
rect 97226 90278 97256 90330
rect 97280 90278 97290 90330
rect 97290 90278 97336 90330
rect 97040 90276 97096 90278
rect 97120 90276 97176 90278
rect 97200 90276 97256 90278
rect 97280 90276 97336 90278
rect 65660 89786 65716 89788
rect 65740 89786 65796 89788
rect 65820 89786 65876 89788
rect 65900 89786 65956 89788
rect 65660 89734 65706 89786
rect 65706 89734 65716 89786
rect 65740 89734 65770 89786
rect 65770 89734 65782 89786
rect 65782 89734 65796 89786
rect 65820 89734 65834 89786
rect 65834 89734 65846 89786
rect 65846 89734 65876 89786
rect 65900 89734 65910 89786
rect 65910 89734 65956 89786
rect 65660 89732 65716 89734
rect 65740 89732 65796 89734
rect 65820 89732 65876 89734
rect 65900 89732 65956 89734
rect 96380 89786 96436 89788
rect 96460 89786 96516 89788
rect 96540 89786 96596 89788
rect 96620 89786 96676 89788
rect 96380 89734 96426 89786
rect 96426 89734 96436 89786
rect 96460 89734 96490 89786
rect 96490 89734 96502 89786
rect 96502 89734 96516 89786
rect 96540 89734 96554 89786
rect 96554 89734 96566 89786
rect 96566 89734 96596 89786
rect 96620 89734 96630 89786
rect 96630 89734 96676 89786
rect 96380 89732 96436 89734
rect 96460 89732 96516 89734
rect 96540 89732 96596 89734
rect 96620 89732 96676 89734
rect 66320 89242 66376 89244
rect 66400 89242 66456 89244
rect 66480 89242 66536 89244
rect 66560 89242 66616 89244
rect 66320 89190 66366 89242
rect 66366 89190 66376 89242
rect 66400 89190 66430 89242
rect 66430 89190 66442 89242
rect 66442 89190 66456 89242
rect 66480 89190 66494 89242
rect 66494 89190 66506 89242
rect 66506 89190 66536 89242
rect 66560 89190 66570 89242
rect 66570 89190 66616 89242
rect 66320 89188 66376 89190
rect 66400 89188 66456 89190
rect 66480 89188 66536 89190
rect 66560 89188 66616 89190
rect 97040 89242 97096 89244
rect 97120 89242 97176 89244
rect 97200 89242 97256 89244
rect 97280 89242 97336 89244
rect 97040 89190 97086 89242
rect 97086 89190 97096 89242
rect 97120 89190 97150 89242
rect 97150 89190 97162 89242
rect 97162 89190 97176 89242
rect 97200 89190 97214 89242
rect 97214 89190 97226 89242
rect 97226 89190 97256 89242
rect 97280 89190 97290 89242
rect 97290 89190 97336 89242
rect 97040 89188 97096 89190
rect 97120 89188 97176 89190
rect 97200 89188 97256 89190
rect 97280 89188 97336 89190
rect 65660 88698 65716 88700
rect 65740 88698 65796 88700
rect 65820 88698 65876 88700
rect 65900 88698 65956 88700
rect 65660 88646 65706 88698
rect 65706 88646 65716 88698
rect 65740 88646 65770 88698
rect 65770 88646 65782 88698
rect 65782 88646 65796 88698
rect 65820 88646 65834 88698
rect 65834 88646 65846 88698
rect 65846 88646 65876 88698
rect 65900 88646 65910 88698
rect 65910 88646 65956 88698
rect 65660 88644 65716 88646
rect 65740 88644 65796 88646
rect 65820 88644 65876 88646
rect 65900 88644 65956 88646
rect 96380 88698 96436 88700
rect 96460 88698 96516 88700
rect 96540 88698 96596 88700
rect 96620 88698 96676 88700
rect 96380 88646 96426 88698
rect 96426 88646 96436 88698
rect 96460 88646 96490 88698
rect 96490 88646 96502 88698
rect 96502 88646 96516 88698
rect 96540 88646 96554 88698
rect 96554 88646 96566 88698
rect 96566 88646 96596 88698
rect 96620 88646 96630 88698
rect 96630 88646 96676 88698
rect 96380 88644 96436 88646
rect 96460 88644 96516 88646
rect 96540 88644 96596 88646
rect 96620 88644 96676 88646
rect 66320 88154 66376 88156
rect 66400 88154 66456 88156
rect 66480 88154 66536 88156
rect 66560 88154 66616 88156
rect 66320 88102 66366 88154
rect 66366 88102 66376 88154
rect 66400 88102 66430 88154
rect 66430 88102 66442 88154
rect 66442 88102 66456 88154
rect 66480 88102 66494 88154
rect 66494 88102 66506 88154
rect 66506 88102 66536 88154
rect 66560 88102 66570 88154
rect 66570 88102 66616 88154
rect 66320 88100 66376 88102
rect 66400 88100 66456 88102
rect 66480 88100 66536 88102
rect 66560 88100 66616 88102
rect 97040 88154 97096 88156
rect 97120 88154 97176 88156
rect 97200 88154 97256 88156
rect 97280 88154 97336 88156
rect 97040 88102 97086 88154
rect 97086 88102 97096 88154
rect 97120 88102 97150 88154
rect 97150 88102 97162 88154
rect 97162 88102 97176 88154
rect 97200 88102 97214 88154
rect 97214 88102 97226 88154
rect 97226 88102 97256 88154
rect 97280 88102 97290 88154
rect 97290 88102 97336 88154
rect 97040 88100 97096 88102
rect 97120 88100 97176 88102
rect 97200 88100 97256 88102
rect 97280 88100 97336 88102
rect 65660 87610 65716 87612
rect 65740 87610 65796 87612
rect 65820 87610 65876 87612
rect 65900 87610 65956 87612
rect 65660 87558 65706 87610
rect 65706 87558 65716 87610
rect 65740 87558 65770 87610
rect 65770 87558 65782 87610
rect 65782 87558 65796 87610
rect 65820 87558 65834 87610
rect 65834 87558 65846 87610
rect 65846 87558 65876 87610
rect 65900 87558 65910 87610
rect 65910 87558 65956 87610
rect 65660 87556 65716 87558
rect 65740 87556 65796 87558
rect 65820 87556 65876 87558
rect 65900 87556 65956 87558
rect 96380 87610 96436 87612
rect 96460 87610 96516 87612
rect 96540 87610 96596 87612
rect 96620 87610 96676 87612
rect 96380 87558 96426 87610
rect 96426 87558 96436 87610
rect 96460 87558 96490 87610
rect 96490 87558 96502 87610
rect 96502 87558 96516 87610
rect 96540 87558 96554 87610
rect 96554 87558 96566 87610
rect 96566 87558 96596 87610
rect 96620 87558 96630 87610
rect 96630 87558 96676 87610
rect 96380 87556 96436 87558
rect 96460 87556 96516 87558
rect 96540 87556 96596 87558
rect 96620 87556 96676 87558
rect 66320 87066 66376 87068
rect 66400 87066 66456 87068
rect 66480 87066 66536 87068
rect 66560 87066 66616 87068
rect 66320 87014 66366 87066
rect 66366 87014 66376 87066
rect 66400 87014 66430 87066
rect 66430 87014 66442 87066
rect 66442 87014 66456 87066
rect 66480 87014 66494 87066
rect 66494 87014 66506 87066
rect 66506 87014 66536 87066
rect 66560 87014 66570 87066
rect 66570 87014 66616 87066
rect 66320 87012 66376 87014
rect 66400 87012 66456 87014
rect 66480 87012 66536 87014
rect 66560 87012 66616 87014
rect 97040 87066 97096 87068
rect 97120 87066 97176 87068
rect 97200 87066 97256 87068
rect 97280 87066 97336 87068
rect 97040 87014 97086 87066
rect 97086 87014 97096 87066
rect 97120 87014 97150 87066
rect 97150 87014 97162 87066
rect 97162 87014 97176 87066
rect 97200 87014 97214 87066
rect 97214 87014 97226 87066
rect 97226 87014 97256 87066
rect 97280 87014 97290 87066
rect 97290 87014 97336 87066
rect 97040 87012 97096 87014
rect 97120 87012 97176 87014
rect 97200 87012 97256 87014
rect 97280 87012 97336 87014
rect 65660 86522 65716 86524
rect 65740 86522 65796 86524
rect 65820 86522 65876 86524
rect 65900 86522 65956 86524
rect 65660 86470 65706 86522
rect 65706 86470 65716 86522
rect 65740 86470 65770 86522
rect 65770 86470 65782 86522
rect 65782 86470 65796 86522
rect 65820 86470 65834 86522
rect 65834 86470 65846 86522
rect 65846 86470 65876 86522
rect 65900 86470 65910 86522
rect 65910 86470 65956 86522
rect 65660 86468 65716 86470
rect 65740 86468 65796 86470
rect 65820 86468 65876 86470
rect 65900 86468 65956 86470
rect 96380 86522 96436 86524
rect 96460 86522 96516 86524
rect 96540 86522 96596 86524
rect 96620 86522 96676 86524
rect 96380 86470 96426 86522
rect 96426 86470 96436 86522
rect 96460 86470 96490 86522
rect 96490 86470 96502 86522
rect 96502 86470 96516 86522
rect 96540 86470 96554 86522
rect 96554 86470 96566 86522
rect 96566 86470 96596 86522
rect 96620 86470 96630 86522
rect 96630 86470 96676 86522
rect 96380 86468 96436 86470
rect 96460 86468 96516 86470
rect 96540 86468 96596 86470
rect 96620 86468 96676 86470
rect 66320 85978 66376 85980
rect 66400 85978 66456 85980
rect 66480 85978 66536 85980
rect 66560 85978 66616 85980
rect 66320 85926 66366 85978
rect 66366 85926 66376 85978
rect 66400 85926 66430 85978
rect 66430 85926 66442 85978
rect 66442 85926 66456 85978
rect 66480 85926 66494 85978
rect 66494 85926 66506 85978
rect 66506 85926 66536 85978
rect 66560 85926 66570 85978
rect 66570 85926 66616 85978
rect 66320 85924 66376 85926
rect 66400 85924 66456 85926
rect 66480 85924 66536 85926
rect 66560 85924 66616 85926
rect 97040 85978 97096 85980
rect 97120 85978 97176 85980
rect 97200 85978 97256 85980
rect 97280 85978 97336 85980
rect 97040 85926 97086 85978
rect 97086 85926 97096 85978
rect 97120 85926 97150 85978
rect 97150 85926 97162 85978
rect 97162 85926 97176 85978
rect 97200 85926 97214 85978
rect 97214 85926 97226 85978
rect 97226 85926 97256 85978
rect 97280 85926 97290 85978
rect 97290 85926 97336 85978
rect 97040 85924 97096 85926
rect 97120 85924 97176 85926
rect 97200 85924 97256 85926
rect 97280 85924 97336 85926
rect 65660 85434 65716 85436
rect 65740 85434 65796 85436
rect 65820 85434 65876 85436
rect 65900 85434 65956 85436
rect 65660 85382 65706 85434
rect 65706 85382 65716 85434
rect 65740 85382 65770 85434
rect 65770 85382 65782 85434
rect 65782 85382 65796 85434
rect 65820 85382 65834 85434
rect 65834 85382 65846 85434
rect 65846 85382 65876 85434
rect 65900 85382 65910 85434
rect 65910 85382 65956 85434
rect 65660 85380 65716 85382
rect 65740 85380 65796 85382
rect 65820 85380 65876 85382
rect 65900 85380 65956 85382
rect 96380 85434 96436 85436
rect 96460 85434 96516 85436
rect 96540 85434 96596 85436
rect 96620 85434 96676 85436
rect 96380 85382 96426 85434
rect 96426 85382 96436 85434
rect 96460 85382 96490 85434
rect 96490 85382 96502 85434
rect 96502 85382 96516 85434
rect 96540 85382 96554 85434
rect 96554 85382 96566 85434
rect 96566 85382 96596 85434
rect 96620 85382 96630 85434
rect 96630 85382 96676 85434
rect 96380 85380 96436 85382
rect 96460 85380 96516 85382
rect 96540 85380 96596 85382
rect 96620 85380 96676 85382
rect 66320 84890 66376 84892
rect 66400 84890 66456 84892
rect 66480 84890 66536 84892
rect 66560 84890 66616 84892
rect 66320 84838 66366 84890
rect 66366 84838 66376 84890
rect 66400 84838 66430 84890
rect 66430 84838 66442 84890
rect 66442 84838 66456 84890
rect 66480 84838 66494 84890
rect 66494 84838 66506 84890
rect 66506 84838 66536 84890
rect 66560 84838 66570 84890
rect 66570 84838 66616 84890
rect 66320 84836 66376 84838
rect 66400 84836 66456 84838
rect 66480 84836 66536 84838
rect 66560 84836 66616 84838
rect 97040 84890 97096 84892
rect 97120 84890 97176 84892
rect 97200 84890 97256 84892
rect 97280 84890 97336 84892
rect 97040 84838 97086 84890
rect 97086 84838 97096 84890
rect 97120 84838 97150 84890
rect 97150 84838 97162 84890
rect 97162 84838 97176 84890
rect 97200 84838 97214 84890
rect 97214 84838 97226 84890
rect 97226 84838 97256 84890
rect 97280 84838 97290 84890
rect 97290 84838 97336 84890
rect 97040 84836 97096 84838
rect 97120 84836 97176 84838
rect 97200 84836 97256 84838
rect 97280 84836 97336 84838
rect 65660 84346 65716 84348
rect 65740 84346 65796 84348
rect 65820 84346 65876 84348
rect 65900 84346 65956 84348
rect 65660 84294 65706 84346
rect 65706 84294 65716 84346
rect 65740 84294 65770 84346
rect 65770 84294 65782 84346
rect 65782 84294 65796 84346
rect 65820 84294 65834 84346
rect 65834 84294 65846 84346
rect 65846 84294 65876 84346
rect 65900 84294 65910 84346
rect 65910 84294 65956 84346
rect 65660 84292 65716 84294
rect 65740 84292 65796 84294
rect 65820 84292 65876 84294
rect 65900 84292 65956 84294
rect 96380 84346 96436 84348
rect 96460 84346 96516 84348
rect 96540 84346 96596 84348
rect 96620 84346 96676 84348
rect 96380 84294 96426 84346
rect 96426 84294 96436 84346
rect 96460 84294 96490 84346
rect 96490 84294 96502 84346
rect 96502 84294 96516 84346
rect 96540 84294 96554 84346
rect 96554 84294 96566 84346
rect 96566 84294 96596 84346
rect 96620 84294 96630 84346
rect 96630 84294 96676 84346
rect 96380 84292 96436 84294
rect 96460 84292 96516 84294
rect 96540 84292 96596 84294
rect 96620 84292 96676 84294
rect 66320 83802 66376 83804
rect 66400 83802 66456 83804
rect 66480 83802 66536 83804
rect 66560 83802 66616 83804
rect 66320 83750 66366 83802
rect 66366 83750 66376 83802
rect 66400 83750 66430 83802
rect 66430 83750 66442 83802
rect 66442 83750 66456 83802
rect 66480 83750 66494 83802
rect 66494 83750 66506 83802
rect 66506 83750 66536 83802
rect 66560 83750 66570 83802
rect 66570 83750 66616 83802
rect 66320 83748 66376 83750
rect 66400 83748 66456 83750
rect 66480 83748 66536 83750
rect 66560 83748 66616 83750
rect 97040 83802 97096 83804
rect 97120 83802 97176 83804
rect 97200 83802 97256 83804
rect 97280 83802 97336 83804
rect 97040 83750 97086 83802
rect 97086 83750 97096 83802
rect 97120 83750 97150 83802
rect 97150 83750 97162 83802
rect 97162 83750 97176 83802
rect 97200 83750 97214 83802
rect 97214 83750 97226 83802
rect 97226 83750 97256 83802
rect 97280 83750 97290 83802
rect 97290 83750 97336 83802
rect 97040 83748 97096 83750
rect 97120 83748 97176 83750
rect 97200 83748 97256 83750
rect 97280 83748 97336 83750
rect 65660 83258 65716 83260
rect 65740 83258 65796 83260
rect 65820 83258 65876 83260
rect 65900 83258 65956 83260
rect 65660 83206 65706 83258
rect 65706 83206 65716 83258
rect 65740 83206 65770 83258
rect 65770 83206 65782 83258
rect 65782 83206 65796 83258
rect 65820 83206 65834 83258
rect 65834 83206 65846 83258
rect 65846 83206 65876 83258
rect 65900 83206 65910 83258
rect 65910 83206 65956 83258
rect 65660 83204 65716 83206
rect 65740 83204 65796 83206
rect 65820 83204 65876 83206
rect 65900 83204 65956 83206
rect 96380 83258 96436 83260
rect 96460 83258 96516 83260
rect 96540 83258 96596 83260
rect 96620 83258 96676 83260
rect 96380 83206 96426 83258
rect 96426 83206 96436 83258
rect 96460 83206 96490 83258
rect 96490 83206 96502 83258
rect 96502 83206 96516 83258
rect 96540 83206 96554 83258
rect 96554 83206 96566 83258
rect 96566 83206 96596 83258
rect 96620 83206 96630 83258
rect 96630 83206 96676 83258
rect 96380 83204 96436 83206
rect 96460 83204 96516 83206
rect 96540 83204 96596 83206
rect 96620 83204 96676 83206
rect 66320 82714 66376 82716
rect 66400 82714 66456 82716
rect 66480 82714 66536 82716
rect 66560 82714 66616 82716
rect 66320 82662 66366 82714
rect 66366 82662 66376 82714
rect 66400 82662 66430 82714
rect 66430 82662 66442 82714
rect 66442 82662 66456 82714
rect 66480 82662 66494 82714
rect 66494 82662 66506 82714
rect 66506 82662 66536 82714
rect 66560 82662 66570 82714
rect 66570 82662 66616 82714
rect 66320 82660 66376 82662
rect 66400 82660 66456 82662
rect 66480 82660 66536 82662
rect 66560 82660 66616 82662
rect 97040 82714 97096 82716
rect 97120 82714 97176 82716
rect 97200 82714 97256 82716
rect 97280 82714 97336 82716
rect 97040 82662 97086 82714
rect 97086 82662 97096 82714
rect 97120 82662 97150 82714
rect 97150 82662 97162 82714
rect 97162 82662 97176 82714
rect 97200 82662 97214 82714
rect 97214 82662 97226 82714
rect 97226 82662 97256 82714
rect 97280 82662 97290 82714
rect 97290 82662 97336 82714
rect 97040 82660 97096 82662
rect 97120 82660 97176 82662
rect 97200 82660 97256 82662
rect 97280 82660 97336 82662
rect 65660 82170 65716 82172
rect 65740 82170 65796 82172
rect 65820 82170 65876 82172
rect 65900 82170 65956 82172
rect 65660 82118 65706 82170
rect 65706 82118 65716 82170
rect 65740 82118 65770 82170
rect 65770 82118 65782 82170
rect 65782 82118 65796 82170
rect 65820 82118 65834 82170
rect 65834 82118 65846 82170
rect 65846 82118 65876 82170
rect 65900 82118 65910 82170
rect 65910 82118 65956 82170
rect 65660 82116 65716 82118
rect 65740 82116 65796 82118
rect 65820 82116 65876 82118
rect 65900 82116 65956 82118
rect 96380 82170 96436 82172
rect 96460 82170 96516 82172
rect 96540 82170 96596 82172
rect 96620 82170 96676 82172
rect 96380 82118 96426 82170
rect 96426 82118 96436 82170
rect 96460 82118 96490 82170
rect 96490 82118 96502 82170
rect 96502 82118 96516 82170
rect 96540 82118 96554 82170
rect 96554 82118 96566 82170
rect 96566 82118 96596 82170
rect 96620 82118 96630 82170
rect 96630 82118 96676 82170
rect 96380 82116 96436 82118
rect 96460 82116 96516 82118
rect 96540 82116 96596 82118
rect 96620 82116 96676 82118
rect 66320 81626 66376 81628
rect 66400 81626 66456 81628
rect 66480 81626 66536 81628
rect 66560 81626 66616 81628
rect 66320 81574 66366 81626
rect 66366 81574 66376 81626
rect 66400 81574 66430 81626
rect 66430 81574 66442 81626
rect 66442 81574 66456 81626
rect 66480 81574 66494 81626
rect 66494 81574 66506 81626
rect 66506 81574 66536 81626
rect 66560 81574 66570 81626
rect 66570 81574 66616 81626
rect 66320 81572 66376 81574
rect 66400 81572 66456 81574
rect 66480 81572 66536 81574
rect 66560 81572 66616 81574
rect 97040 81626 97096 81628
rect 97120 81626 97176 81628
rect 97200 81626 97256 81628
rect 97280 81626 97336 81628
rect 97040 81574 97086 81626
rect 97086 81574 97096 81626
rect 97120 81574 97150 81626
rect 97150 81574 97162 81626
rect 97162 81574 97176 81626
rect 97200 81574 97214 81626
rect 97214 81574 97226 81626
rect 97226 81574 97256 81626
rect 97280 81574 97290 81626
rect 97290 81574 97336 81626
rect 97040 81572 97096 81574
rect 97120 81572 97176 81574
rect 97200 81572 97256 81574
rect 97280 81572 97336 81574
rect 65660 81082 65716 81084
rect 65740 81082 65796 81084
rect 65820 81082 65876 81084
rect 65900 81082 65956 81084
rect 65660 81030 65706 81082
rect 65706 81030 65716 81082
rect 65740 81030 65770 81082
rect 65770 81030 65782 81082
rect 65782 81030 65796 81082
rect 65820 81030 65834 81082
rect 65834 81030 65846 81082
rect 65846 81030 65876 81082
rect 65900 81030 65910 81082
rect 65910 81030 65956 81082
rect 65660 81028 65716 81030
rect 65740 81028 65796 81030
rect 65820 81028 65876 81030
rect 65900 81028 65956 81030
rect 96380 81082 96436 81084
rect 96460 81082 96516 81084
rect 96540 81082 96596 81084
rect 96620 81082 96676 81084
rect 96380 81030 96426 81082
rect 96426 81030 96436 81082
rect 96460 81030 96490 81082
rect 96490 81030 96502 81082
rect 96502 81030 96516 81082
rect 96540 81030 96554 81082
rect 96554 81030 96566 81082
rect 96566 81030 96596 81082
rect 96620 81030 96630 81082
rect 96630 81030 96676 81082
rect 96380 81028 96436 81030
rect 96460 81028 96516 81030
rect 96540 81028 96596 81030
rect 96620 81028 96676 81030
rect 66320 80538 66376 80540
rect 66400 80538 66456 80540
rect 66480 80538 66536 80540
rect 66560 80538 66616 80540
rect 66320 80486 66366 80538
rect 66366 80486 66376 80538
rect 66400 80486 66430 80538
rect 66430 80486 66442 80538
rect 66442 80486 66456 80538
rect 66480 80486 66494 80538
rect 66494 80486 66506 80538
rect 66506 80486 66536 80538
rect 66560 80486 66570 80538
rect 66570 80486 66616 80538
rect 66320 80484 66376 80486
rect 66400 80484 66456 80486
rect 66480 80484 66536 80486
rect 66560 80484 66616 80486
rect 97040 80538 97096 80540
rect 97120 80538 97176 80540
rect 97200 80538 97256 80540
rect 97280 80538 97336 80540
rect 97040 80486 97086 80538
rect 97086 80486 97096 80538
rect 97120 80486 97150 80538
rect 97150 80486 97162 80538
rect 97162 80486 97176 80538
rect 97200 80486 97214 80538
rect 97214 80486 97226 80538
rect 97226 80486 97256 80538
rect 97280 80486 97290 80538
rect 97290 80486 97336 80538
rect 97040 80484 97096 80486
rect 97120 80484 97176 80486
rect 97200 80484 97256 80486
rect 97280 80484 97336 80486
rect 65660 79994 65716 79996
rect 65740 79994 65796 79996
rect 65820 79994 65876 79996
rect 65900 79994 65956 79996
rect 65660 79942 65706 79994
rect 65706 79942 65716 79994
rect 65740 79942 65770 79994
rect 65770 79942 65782 79994
rect 65782 79942 65796 79994
rect 65820 79942 65834 79994
rect 65834 79942 65846 79994
rect 65846 79942 65876 79994
rect 65900 79942 65910 79994
rect 65910 79942 65956 79994
rect 65660 79940 65716 79942
rect 65740 79940 65796 79942
rect 65820 79940 65876 79942
rect 65900 79940 65956 79942
rect 96380 79994 96436 79996
rect 96460 79994 96516 79996
rect 96540 79994 96596 79996
rect 96620 79994 96676 79996
rect 96380 79942 96426 79994
rect 96426 79942 96436 79994
rect 96460 79942 96490 79994
rect 96490 79942 96502 79994
rect 96502 79942 96516 79994
rect 96540 79942 96554 79994
rect 96554 79942 96566 79994
rect 96566 79942 96596 79994
rect 96620 79942 96630 79994
rect 96630 79942 96676 79994
rect 96380 79940 96436 79942
rect 96460 79940 96516 79942
rect 96540 79940 96596 79942
rect 96620 79940 96676 79942
rect 66320 79450 66376 79452
rect 66400 79450 66456 79452
rect 66480 79450 66536 79452
rect 66560 79450 66616 79452
rect 66320 79398 66366 79450
rect 66366 79398 66376 79450
rect 66400 79398 66430 79450
rect 66430 79398 66442 79450
rect 66442 79398 66456 79450
rect 66480 79398 66494 79450
rect 66494 79398 66506 79450
rect 66506 79398 66536 79450
rect 66560 79398 66570 79450
rect 66570 79398 66616 79450
rect 66320 79396 66376 79398
rect 66400 79396 66456 79398
rect 66480 79396 66536 79398
rect 66560 79396 66616 79398
rect 97040 79450 97096 79452
rect 97120 79450 97176 79452
rect 97200 79450 97256 79452
rect 97280 79450 97336 79452
rect 97040 79398 97086 79450
rect 97086 79398 97096 79450
rect 97120 79398 97150 79450
rect 97150 79398 97162 79450
rect 97162 79398 97176 79450
rect 97200 79398 97214 79450
rect 97214 79398 97226 79450
rect 97226 79398 97256 79450
rect 97280 79398 97290 79450
rect 97290 79398 97336 79450
rect 97040 79396 97096 79398
rect 97120 79396 97176 79398
rect 97200 79396 97256 79398
rect 97280 79396 97336 79398
rect 65660 78906 65716 78908
rect 65740 78906 65796 78908
rect 65820 78906 65876 78908
rect 65900 78906 65956 78908
rect 65660 78854 65706 78906
rect 65706 78854 65716 78906
rect 65740 78854 65770 78906
rect 65770 78854 65782 78906
rect 65782 78854 65796 78906
rect 65820 78854 65834 78906
rect 65834 78854 65846 78906
rect 65846 78854 65876 78906
rect 65900 78854 65910 78906
rect 65910 78854 65956 78906
rect 65660 78852 65716 78854
rect 65740 78852 65796 78854
rect 65820 78852 65876 78854
rect 65900 78852 65956 78854
rect 96380 78906 96436 78908
rect 96460 78906 96516 78908
rect 96540 78906 96596 78908
rect 96620 78906 96676 78908
rect 96380 78854 96426 78906
rect 96426 78854 96436 78906
rect 96460 78854 96490 78906
rect 96490 78854 96502 78906
rect 96502 78854 96516 78906
rect 96540 78854 96554 78906
rect 96554 78854 96566 78906
rect 96566 78854 96596 78906
rect 96620 78854 96630 78906
rect 96630 78854 96676 78906
rect 96380 78852 96436 78854
rect 96460 78852 96516 78854
rect 96540 78852 96596 78854
rect 96620 78852 96676 78854
rect 66320 78362 66376 78364
rect 66400 78362 66456 78364
rect 66480 78362 66536 78364
rect 66560 78362 66616 78364
rect 66320 78310 66366 78362
rect 66366 78310 66376 78362
rect 66400 78310 66430 78362
rect 66430 78310 66442 78362
rect 66442 78310 66456 78362
rect 66480 78310 66494 78362
rect 66494 78310 66506 78362
rect 66506 78310 66536 78362
rect 66560 78310 66570 78362
rect 66570 78310 66616 78362
rect 66320 78308 66376 78310
rect 66400 78308 66456 78310
rect 66480 78308 66536 78310
rect 66560 78308 66616 78310
rect 97040 78362 97096 78364
rect 97120 78362 97176 78364
rect 97200 78362 97256 78364
rect 97280 78362 97336 78364
rect 97040 78310 97086 78362
rect 97086 78310 97096 78362
rect 97120 78310 97150 78362
rect 97150 78310 97162 78362
rect 97162 78310 97176 78362
rect 97200 78310 97214 78362
rect 97214 78310 97226 78362
rect 97226 78310 97256 78362
rect 97280 78310 97290 78362
rect 97290 78310 97336 78362
rect 97040 78308 97096 78310
rect 97120 78308 97176 78310
rect 97200 78308 97256 78310
rect 97280 78308 97336 78310
rect 65660 77818 65716 77820
rect 65740 77818 65796 77820
rect 65820 77818 65876 77820
rect 65900 77818 65956 77820
rect 65660 77766 65706 77818
rect 65706 77766 65716 77818
rect 65740 77766 65770 77818
rect 65770 77766 65782 77818
rect 65782 77766 65796 77818
rect 65820 77766 65834 77818
rect 65834 77766 65846 77818
rect 65846 77766 65876 77818
rect 65900 77766 65910 77818
rect 65910 77766 65956 77818
rect 65660 77764 65716 77766
rect 65740 77764 65796 77766
rect 65820 77764 65876 77766
rect 65900 77764 65956 77766
rect 96380 77818 96436 77820
rect 96460 77818 96516 77820
rect 96540 77818 96596 77820
rect 96620 77818 96676 77820
rect 96380 77766 96426 77818
rect 96426 77766 96436 77818
rect 96460 77766 96490 77818
rect 96490 77766 96502 77818
rect 96502 77766 96516 77818
rect 96540 77766 96554 77818
rect 96554 77766 96566 77818
rect 96566 77766 96596 77818
rect 96620 77766 96630 77818
rect 96630 77766 96676 77818
rect 96380 77764 96436 77766
rect 96460 77764 96516 77766
rect 96540 77764 96596 77766
rect 96620 77764 96676 77766
rect 53286 75792 53342 75848
rect 55586 74568 55642 74624
rect 66320 77274 66376 77276
rect 66400 77274 66456 77276
rect 66480 77274 66536 77276
rect 66560 77274 66616 77276
rect 66320 77222 66366 77274
rect 66366 77222 66376 77274
rect 66400 77222 66430 77274
rect 66430 77222 66442 77274
rect 66442 77222 66456 77274
rect 66480 77222 66494 77274
rect 66494 77222 66506 77274
rect 66506 77222 66536 77274
rect 66560 77222 66570 77274
rect 66570 77222 66616 77274
rect 66320 77220 66376 77222
rect 66400 77220 66456 77222
rect 66480 77220 66536 77222
rect 66560 77220 66616 77222
rect 97040 77274 97096 77276
rect 97120 77274 97176 77276
rect 97200 77274 97256 77276
rect 97280 77274 97336 77276
rect 97040 77222 97086 77274
rect 97086 77222 97096 77274
rect 97120 77222 97150 77274
rect 97150 77222 97162 77274
rect 97162 77222 97176 77274
rect 97200 77222 97214 77274
rect 97214 77222 97226 77274
rect 97226 77222 97256 77274
rect 97280 77222 97290 77274
rect 97290 77222 97336 77274
rect 97040 77220 97096 77222
rect 97120 77220 97176 77222
rect 97200 77220 97256 77222
rect 97280 77220 97336 77222
rect 65660 76730 65716 76732
rect 65740 76730 65796 76732
rect 65820 76730 65876 76732
rect 65900 76730 65956 76732
rect 65660 76678 65706 76730
rect 65706 76678 65716 76730
rect 65740 76678 65770 76730
rect 65770 76678 65782 76730
rect 65782 76678 65796 76730
rect 65820 76678 65834 76730
rect 65834 76678 65846 76730
rect 65846 76678 65876 76730
rect 65900 76678 65910 76730
rect 65910 76678 65956 76730
rect 65660 76676 65716 76678
rect 65740 76676 65796 76678
rect 65820 76676 65876 76678
rect 65900 76676 65956 76678
rect 96380 76730 96436 76732
rect 96460 76730 96516 76732
rect 96540 76730 96596 76732
rect 96620 76730 96676 76732
rect 96380 76678 96426 76730
rect 96426 76678 96436 76730
rect 96460 76678 96490 76730
rect 96490 76678 96502 76730
rect 96502 76678 96516 76730
rect 96540 76678 96554 76730
rect 96554 76678 96566 76730
rect 96566 76678 96596 76730
rect 96620 76678 96630 76730
rect 96630 76678 96676 76730
rect 96380 76676 96436 76678
rect 96460 76676 96516 76678
rect 96540 76676 96596 76678
rect 96620 76676 96676 76678
rect 66320 76186 66376 76188
rect 66400 76186 66456 76188
rect 66480 76186 66536 76188
rect 66560 76186 66616 76188
rect 66320 76134 66366 76186
rect 66366 76134 66376 76186
rect 66400 76134 66430 76186
rect 66430 76134 66442 76186
rect 66442 76134 66456 76186
rect 66480 76134 66494 76186
rect 66494 76134 66506 76186
rect 66506 76134 66536 76186
rect 66560 76134 66570 76186
rect 66570 76134 66616 76186
rect 66320 76132 66376 76134
rect 66400 76132 66456 76134
rect 66480 76132 66536 76134
rect 66560 76132 66616 76134
rect 97040 76186 97096 76188
rect 97120 76186 97176 76188
rect 97200 76186 97256 76188
rect 97280 76186 97336 76188
rect 97040 76134 97086 76186
rect 97086 76134 97096 76186
rect 97120 76134 97150 76186
rect 97150 76134 97162 76186
rect 97162 76134 97176 76186
rect 97200 76134 97214 76186
rect 97214 76134 97226 76186
rect 97226 76134 97256 76186
rect 97280 76134 97290 76186
rect 97290 76134 97336 76186
rect 97040 76132 97096 76134
rect 97120 76132 97176 76134
rect 97200 76132 97256 76134
rect 97280 76132 97336 76134
rect 65660 75642 65716 75644
rect 65740 75642 65796 75644
rect 65820 75642 65876 75644
rect 65900 75642 65956 75644
rect 65660 75590 65706 75642
rect 65706 75590 65716 75642
rect 65740 75590 65770 75642
rect 65770 75590 65782 75642
rect 65782 75590 65796 75642
rect 65820 75590 65834 75642
rect 65834 75590 65846 75642
rect 65846 75590 65876 75642
rect 65900 75590 65910 75642
rect 65910 75590 65956 75642
rect 65660 75588 65716 75590
rect 65740 75588 65796 75590
rect 65820 75588 65876 75590
rect 65900 75588 65956 75590
rect 96380 75642 96436 75644
rect 96460 75642 96516 75644
rect 96540 75642 96596 75644
rect 96620 75642 96676 75644
rect 96380 75590 96426 75642
rect 96426 75590 96436 75642
rect 96460 75590 96490 75642
rect 96490 75590 96502 75642
rect 96502 75590 96516 75642
rect 96540 75590 96554 75642
rect 96554 75590 96566 75642
rect 96566 75590 96596 75642
rect 96620 75590 96630 75642
rect 96630 75590 96676 75642
rect 96380 75588 96436 75590
rect 96460 75588 96516 75590
rect 96540 75588 96596 75590
rect 96620 75588 96676 75590
rect 66320 75098 66376 75100
rect 66400 75098 66456 75100
rect 66480 75098 66536 75100
rect 66560 75098 66616 75100
rect 66320 75046 66366 75098
rect 66366 75046 66376 75098
rect 66400 75046 66430 75098
rect 66430 75046 66442 75098
rect 66442 75046 66456 75098
rect 66480 75046 66494 75098
rect 66494 75046 66506 75098
rect 66506 75046 66536 75098
rect 66560 75046 66570 75098
rect 66570 75046 66616 75098
rect 66320 75044 66376 75046
rect 66400 75044 66456 75046
rect 66480 75044 66536 75046
rect 66560 75044 66616 75046
rect 97040 75098 97096 75100
rect 97120 75098 97176 75100
rect 97200 75098 97256 75100
rect 97280 75098 97336 75100
rect 97040 75046 97086 75098
rect 97086 75046 97096 75098
rect 97120 75046 97150 75098
rect 97150 75046 97162 75098
rect 97162 75046 97176 75098
rect 97200 75046 97214 75098
rect 97214 75046 97226 75098
rect 97226 75046 97256 75098
rect 97280 75046 97290 75098
rect 97290 75046 97336 75098
rect 97040 75044 97096 75046
rect 97120 75044 97176 75046
rect 97200 75044 97256 75046
rect 97280 75044 97336 75046
rect 65660 74554 65716 74556
rect 65740 74554 65796 74556
rect 65820 74554 65876 74556
rect 65900 74554 65956 74556
rect 65660 74502 65706 74554
rect 65706 74502 65716 74554
rect 65740 74502 65770 74554
rect 65770 74502 65782 74554
rect 65782 74502 65796 74554
rect 65820 74502 65834 74554
rect 65834 74502 65846 74554
rect 65846 74502 65876 74554
rect 65900 74502 65910 74554
rect 65910 74502 65956 74554
rect 65660 74500 65716 74502
rect 65740 74500 65796 74502
rect 65820 74500 65876 74502
rect 65900 74500 65956 74502
rect 66320 74010 66376 74012
rect 66400 74010 66456 74012
rect 66480 74010 66536 74012
rect 66560 74010 66616 74012
rect 66320 73958 66366 74010
rect 66366 73958 66376 74010
rect 66400 73958 66430 74010
rect 66430 73958 66442 74010
rect 66442 73958 66456 74010
rect 66480 73958 66494 74010
rect 66494 73958 66506 74010
rect 66506 73958 66536 74010
rect 66560 73958 66570 74010
rect 66570 73958 66616 74010
rect 66320 73956 66376 73958
rect 66400 73956 66456 73958
rect 66480 73956 66536 73958
rect 66560 73956 66616 73958
rect 57518 73888 57574 73944
rect 65660 73466 65716 73468
rect 65740 73466 65796 73468
rect 65820 73466 65876 73468
rect 65900 73466 65956 73468
rect 65660 73414 65706 73466
rect 65706 73414 65716 73466
rect 65740 73414 65770 73466
rect 65770 73414 65782 73466
rect 65782 73414 65796 73466
rect 65820 73414 65834 73466
rect 65834 73414 65846 73466
rect 65846 73414 65876 73466
rect 65900 73414 65910 73466
rect 65910 73414 65956 73466
rect 65660 73412 65716 73414
rect 65740 73412 65796 73414
rect 65820 73412 65876 73414
rect 65900 73412 65956 73414
rect 66320 72922 66376 72924
rect 66400 72922 66456 72924
rect 66480 72922 66536 72924
rect 66560 72922 66616 72924
rect 66320 72870 66366 72922
rect 66366 72870 66376 72922
rect 66400 72870 66430 72922
rect 66430 72870 66442 72922
rect 66442 72870 66456 72922
rect 66480 72870 66494 72922
rect 66494 72870 66506 72922
rect 66506 72870 66536 72922
rect 66560 72870 66570 72922
rect 66570 72870 66616 72922
rect 66320 72868 66376 72870
rect 66400 72868 66456 72870
rect 66480 72868 66536 72870
rect 66560 72868 66616 72870
rect 65660 72378 65716 72380
rect 65740 72378 65796 72380
rect 65820 72378 65876 72380
rect 65900 72378 65956 72380
rect 65660 72326 65706 72378
rect 65706 72326 65716 72378
rect 65740 72326 65770 72378
rect 65770 72326 65782 72378
rect 65782 72326 65796 72378
rect 65820 72326 65834 72378
rect 65834 72326 65846 72378
rect 65846 72326 65876 72378
rect 65900 72326 65910 72378
rect 65910 72326 65956 72378
rect 65660 72324 65716 72326
rect 65740 72324 65796 72326
rect 65820 72324 65876 72326
rect 65900 72324 65956 72326
rect 51262 71848 51318 71904
rect 66320 71834 66376 71836
rect 66400 71834 66456 71836
rect 66480 71834 66536 71836
rect 66560 71834 66616 71836
rect 66320 71782 66366 71834
rect 66366 71782 66376 71834
rect 66400 71782 66430 71834
rect 66430 71782 66442 71834
rect 66442 71782 66456 71834
rect 66480 71782 66494 71834
rect 66494 71782 66506 71834
rect 66506 71782 66536 71834
rect 66560 71782 66570 71834
rect 66570 71782 66616 71834
rect 66320 71780 66376 71782
rect 66400 71780 66456 71782
rect 66480 71780 66536 71782
rect 66560 71780 66616 71782
rect 65660 71290 65716 71292
rect 65740 71290 65796 71292
rect 65820 71290 65876 71292
rect 65900 71290 65956 71292
rect 65660 71238 65706 71290
rect 65706 71238 65716 71290
rect 65740 71238 65770 71290
rect 65770 71238 65782 71290
rect 65782 71238 65796 71290
rect 65820 71238 65834 71290
rect 65834 71238 65846 71290
rect 65846 71238 65876 71290
rect 65900 71238 65910 71290
rect 65910 71238 65956 71290
rect 65660 71236 65716 71238
rect 65740 71236 65796 71238
rect 65820 71236 65876 71238
rect 65900 71236 65956 71238
rect 66320 70746 66376 70748
rect 66400 70746 66456 70748
rect 66480 70746 66536 70748
rect 66560 70746 66616 70748
rect 66320 70694 66366 70746
rect 66366 70694 66376 70746
rect 66400 70694 66430 70746
rect 66430 70694 66442 70746
rect 66442 70694 66456 70746
rect 66480 70694 66494 70746
rect 66494 70694 66506 70746
rect 66506 70694 66536 70746
rect 66560 70694 66570 70746
rect 66570 70694 66616 70746
rect 66320 70692 66376 70694
rect 66400 70692 66456 70694
rect 66480 70692 66536 70694
rect 66560 70692 66616 70694
rect 65660 70202 65716 70204
rect 65740 70202 65796 70204
rect 65820 70202 65876 70204
rect 65900 70202 65956 70204
rect 65660 70150 65706 70202
rect 65706 70150 65716 70202
rect 65740 70150 65770 70202
rect 65770 70150 65782 70202
rect 65782 70150 65796 70202
rect 65820 70150 65834 70202
rect 65834 70150 65846 70202
rect 65846 70150 65876 70202
rect 65900 70150 65910 70202
rect 65910 70150 65956 70202
rect 65660 70148 65716 70150
rect 65740 70148 65796 70150
rect 65820 70148 65876 70150
rect 65900 70148 65956 70150
rect 66320 69658 66376 69660
rect 66400 69658 66456 69660
rect 66480 69658 66536 69660
rect 66560 69658 66616 69660
rect 66320 69606 66366 69658
rect 66366 69606 66376 69658
rect 66400 69606 66430 69658
rect 66430 69606 66442 69658
rect 66442 69606 66456 69658
rect 66480 69606 66494 69658
rect 66494 69606 66506 69658
rect 66506 69606 66536 69658
rect 66560 69606 66570 69658
rect 66570 69606 66616 69658
rect 66320 69604 66376 69606
rect 66400 69604 66456 69606
rect 66480 69604 66536 69606
rect 66560 69604 66616 69606
rect 65660 69114 65716 69116
rect 65740 69114 65796 69116
rect 65820 69114 65876 69116
rect 65900 69114 65956 69116
rect 65660 69062 65706 69114
rect 65706 69062 65716 69114
rect 65740 69062 65770 69114
rect 65770 69062 65782 69114
rect 65782 69062 65796 69114
rect 65820 69062 65834 69114
rect 65834 69062 65846 69114
rect 65846 69062 65876 69114
rect 65900 69062 65910 69114
rect 65910 69062 65956 69114
rect 65660 69060 65716 69062
rect 65740 69060 65796 69062
rect 65820 69060 65876 69062
rect 65900 69060 65956 69062
rect 66320 68570 66376 68572
rect 66400 68570 66456 68572
rect 66480 68570 66536 68572
rect 66560 68570 66616 68572
rect 66320 68518 66366 68570
rect 66366 68518 66376 68570
rect 66400 68518 66430 68570
rect 66430 68518 66442 68570
rect 66442 68518 66456 68570
rect 66480 68518 66494 68570
rect 66494 68518 66506 68570
rect 66506 68518 66536 68570
rect 66560 68518 66570 68570
rect 66570 68518 66616 68570
rect 66320 68516 66376 68518
rect 66400 68516 66456 68518
rect 66480 68516 66536 68518
rect 66560 68516 66616 68518
rect 65660 68026 65716 68028
rect 65740 68026 65796 68028
rect 65820 68026 65876 68028
rect 65900 68026 65956 68028
rect 65660 67974 65706 68026
rect 65706 67974 65716 68026
rect 65740 67974 65770 68026
rect 65770 67974 65782 68026
rect 65782 67974 65796 68026
rect 65820 67974 65834 68026
rect 65834 67974 65846 68026
rect 65846 67974 65876 68026
rect 65900 67974 65910 68026
rect 65910 67974 65956 68026
rect 65660 67972 65716 67974
rect 65740 67972 65796 67974
rect 65820 67972 65876 67974
rect 65900 67972 65956 67974
rect 66320 67482 66376 67484
rect 66400 67482 66456 67484
rect 66480 67482 66536 67484
rect 66560 67482 66616 67484
rect 66320 67430 66366 67482
rect 66366 67430 66376 67482
rect 66400 67430 66430 67482
rect 66430 67430 66442 67482
rect 66442 67430 66456 67482
rect 66480 67430 66494 67482
rect 66494 67430 66506 67482
rect 66506 67430 66536 67482
rect 66560 67430 66570 67482
rect 66570 67430 66616 67482
rect 66320 67428 66376 67430
rect 66400 67428 66456 67430
rect 66480 67428 66536 67430
rect 66560 67428 66616 67430
rect 65660 66938 65716 66940
rect 65740 66938 65796 66940
rect 65820 66938 65876 66940
rect 65900 66938 65956 66940
rect 65660 66886 65706 66938
rect 65706 66886 65716 66938
rect 65740 66886 65770 66938
rect 65770 66886 65782 66938
rect 65782 66886 65796 66938
rect 65820 66886 65834 66938
rect 65834 66886 65846 66938
rect 65846 66886 65876 66938
rect 65900 66886 65910 66938
rect 65910 66886 65956 66938
rect 65660 66884 65716 66886
rect 65740 66884 65796 66886
rect 65820 66884 65876 66886
rect 65900 66884 65956 66886
rect 66320 66394 66376 66396
rect 66400 66394 66456 66396
rect 66480 66394 66536 66396
rect 66560 66394 66616 66396
rect 66320 66342 66366 66394
rect 66366 66342 66376 66394
rect 66400 66342 66430 66394
rect 66430 66342 66442 66394
rect 66442 66342 66456 66394
rect 66480 66342 66494 66394
rect 66494 66342 66506 66394
rect 66506 66342 66536 66394
rect 66560 66342 66570 66394
rect 66570 66342 66616 66394
rect 66320 66340 66376 66342
rect 66400 66340 66456 66342
rect 66480 66340 66536 66342
rect 66560 66340 66616 66342
rect 65660 65850 65716 65852
rect 65740 65850 65796 65852
rect 65820 65850 65876 65852
rect 65900 65850 65956 65852
rect 65660 65798 65706 65850
rect 65706 65798 65716 65850
rect 65740 65798 65770 65850
rect 65770 65798 65782 65850
rect 65782 65798 65796 65850
rect 65820 65798 65834 65850
rect 65834 65798 65846 65850
rect 65846 65798 65876 65850
rect 65900 65798 65910 65850
rect 65910 65798 65956 65850
rect 65660 65796 65716 65798
rect 65740 65796 65796 65798
rect 65820 65796 65876 65798
rect 65900 65796 65956 65798
rect 66320 65306 66376 65308
rect 66400 65306 66456 65308
rect 66480 65306 66536 65308
rect 66560 65306 66616 65308
rect 66320 65254 66366 65306
rect 66366 65254 66376 65306
rect 66400 65254 66430 65306
rect 66430 65254 66442 65306
rect 66442 65254 66456 65306
rect 66480 65254 66494 65306
rect 66494 65254 66506 65306
rect 66506 65254 66536 65306
rect 66560 65254 66570 65306
rect 66570 65254 66616 65306
rect 66320 65252 66376 65254
rect 66400 65252 66456 65254
rect 66480 65252 66536 65254
rect 66560 65252 66616 65254
rect 65660 64762 65716 64764
rect 65740 64762 65796 64764
rect 65820 64762 65876 64764
rect 65900 64762 65956 64764
rect 65660 64710 65706 64762
rect 65706 64710 65716 64762
rect 65740 64710 65770 64762
rect 65770 64710 65782 64762
rect 65782 64710 65796 64762
rect 65820 64710 65834 64762
rect 65834 64710 65846 64762
rect 65846 64710 65876 64762
rect 65900 64710 65910 64762
rect 65910 64710 65956 64762
rect 65660 64708 65716 64710
rect 65740 64708 65796 64710
rect 65820 64708 65876 64710
rect 65900 64708 65956 64710
rect 66320 64218 66376 64220
rect 66400 64218 66456 64220
rect 66480 64218 66536 64220
rect 66560 64218 66616 64220
rect 66320 64166 66366 64218
rect 66366 64166 66376 64218
rect 66400 64166 66430 64218
rect 66430 64166 66442 64218
rect 66442 64166 66456 64218
rect 66480 64166 66494 64218
rect 66494 64166 66506 64218
rect 66506 64166 66536 64218
rect 66560 64166 66570 64218
rect 66570 64166 66616 64218
rect 66320 64164 66376 64166
rect 66400 64164 66456 64166
rect 66480 64164 66536 64166
rect 66560 64164 66616 64166
rect 65660 63674 65716 63676
rect 65740 63674 65796 63676
rect 65820 63674 65876 63676
rect 65900 63674 65956 63676
rect 65660 63622 65706 63674
rect 65706 63622 65716 63674
rect 65740 63622 65770 63674
rect 65770 63622 65782 63674
rect 65782 63622 65796 63674
rect 65820 63622 65834 63674
rect 65834 63622 65846 63674
rect 65846 63622 65876 63674
rect 65900 63622 65910 63674
rect 65910 63622 65956 63674
rect 65660 63620 65716 63622
rect 65740 63620 65796 63622
rect 65820 63620 65876 63622
rect 65900 63620 65956 63622
rect 66320 63130 66376 63132
rect 66400 63130 66456 63132
rect 66480 63130 66536 63132
rect 66560 63130 66616 63132
rect 66320 63078 66366 63130
rect 66366 63078 66376 63130
rect 66400 63078 66430 63130
rect 66430 63078 66442 63130
rect 66442 63078 66456 63130
rect 66480 63078 66494 63130
rect 66494 63078 66506 63130
rect 66506 63078 66536 63130
rect 66560 63078 66570 63130
rect 66570 63078 66616 63130
rect 66320 63076 66376 63078
rect 66400 63076 66456 63078
rect 66480 63076 66536 63078
rect 66560 63076 66616 63078
rect 65660 62586 65716 62588
rect 65740 62586 65796 62588
rect 65820 62586 65876 62588
rect 65900 62586 65956 62588
rect 65660 62534 65706 62586
rect 65706 62534 65716 62586
rect 65740 62534 65770 62586
rect 65770 62534 65782 62586
rect 65782 62534 65796 62586
rect 65820 62534 65834 62586
rect 65834 62534 65846 62586
rect 65846 62534 65876 62586
rect 65900 62534 65910 62586
rect 65910 62534 65956 62586
rect 65660 62532 65716 62534
rect 65740 62532 65796 62534
rect 65820 62532 65876 62534
rect 65900 62532 65956 62534
rect 66320 62042 66376 62044
rect 66400 62042 66456 62044
rect 66480 62042 66536 62044
rect 66560 62042 66616 62044
rect 66320 61990 66366 62042
rect 66366 61990 66376 62042
rect 66400 61990 66430 62042
rect 66430 61990 66442 62042
rect 66442 61990 66456 62042
rect 66480 61990 66494 62042
rect 66494 61990 66506 62042
rect 66506 61990 66536 62042
rect 66560 61990 66570 62042
rect 66570 61990 66616 62042
rect 66320 61988 66376 61990
rect 66400 61988 66456 61990
rect 66480 61988 66536 61990
rect 66560 61988 66616 61990
rect 65660 61498 65716 61500
rect 65740 61498 65796 61500
rect 65820 61498 65876 61500
rect 65900 61498 65956 61500
rect 65660 61446 65706 61498
rect 65706 61446 65716 61498
rect 65740 61446 65770 61498
rect 65770 61446 65782 61498
rect 65782 61446 65796 61498
rect 65820 61446 65834 61498
rect 65834 61446 65846 61498
rect 65846 61446 65876 61498
rect 65900 61446 65910 61498
rect 65910 61446 65956 61498
rect 65660 61444 65716 61446
rect 65740 61444 65796 61446
rect 65820 61444 65876 61446
rect 65900 61444 65956 61446
rect 66320 60954 66376 60956
rect 66400 60954 66456 60956
rect 66480 60954 66536 60956
rect 66560 60954 66616 60956
rect 66320 60902 66366 60954
rect 66366 60902 66376 60954
rect 66400 60902 66430 60954
rect 66430 60902 66442 60954
rect 66442 60902 66456 60954
rect 66480 60902 66494 60954
rect 66494 60902 66506 60954
rect 66506 60902 66536 60954
rect 66560 60902 66570 60954
rect 66570 60902 66616 60954
rect 66320 60900 66376 60902
rect 66400 60900 66456 60902
rect 66480 60900 66536 60902
rect 66560 60900 66616 60902
rect 34940 60410 34996 60412
rect 35020 60410 35076 60412
rect 35100 60410 35156 60412
rect 35180 60410 35236 60412
rect 34940 60358 34986 60410
rect 34986 60358 34996 60410
rect 35020 60358 35050 60410
rect 35050 60358 35062 60410
rect 35062 60358 35076 60410
rect 35100 60358 35114 60410
rect 35114 60358 35126 60410
rect 35126 60358 35156 60410
rect 35180 60358 35190 60410
rect 35190 60358 35236 60410
rect 34940 60356 34996 60358
rect 35020 60356 35076 60358
rect 35100 60356 35156 60358
rect 35180 60356 35236 60358
rect 65660 60410 65716 60412
rect 65740 60410 65796 60412
rect 65820 60410 65876 60412
rect 65900 60410 65956 60412
rect 65660 60358 65706 60410
rect 65706 60358 65716 60410
rect 65740 60358 65770 60410
rect 65770 60358 65782 60410
rect 65782 60358 65796 60410
rect 65820 60358 65834 60410
rect 65834 60358 65846 60410
rect 65846 60358 65876 60410
rect 65900 60358 65910 60410
rect 65910 60358 65956 60410
rect 65660 60356 65716 60358
rect 65740 60356 65796 60358
rect 65820 60356 65876 60358
rect 65900 60356 65956 60358
rect 35600 59866 35656 59868
rect 35680 59866 35736 59868
rect 35760 59866 35816 59868
rect 35840 59866 35896 59868
rect 35600 59814 35646 59866
rect 35646 59814 35656 59866
rect 35680 59814 35710 59866
rect 35710 59814 35722 59866
rect 35722 59814 35736 59866
rect 35760 59814 35774 59866
rect 35774 59814 35786 59866
rect 35786 59814 35816 59866
rect 35840 59814 35850 59866
rect 35850 59814 35896 59866
rect 35600 59812 35656 59814
rect 35680 59812 35736 59814
rect 35760 59812 35816 59814
rect 35840 59812 35896 59814
rect 66320 59866 66376 59868
rect 66400 59866 66456 59868
rect 66480 59866 66536 59868
rect 66560 59866 66616 59868
rect 66320 59814 66366 59866
rect 66366 59814 66376 59866
rect 66400 59814 66430 59866
rect 66430 59814 66442 59866
rect 66442 59814 66456 59866
rect 66480 59814 66494 59866
rect 66494 59814 66506 59866
rect 66506 59814 66536 59866
rect 66560 59814 66570 59866
rect 66570 59814 66616 59866
rect 66320 59812 66376 59814
rect 66400 59812 66456 59814
rect 66480 59812 66536 59814
rect 66560 59812 66616 59814
rect 77114 60696 77170 60752
rect 71778 58792 71834 58848
rect 96380 74554 96436 74556
rect 96460 74554 96516 74556
rect 96540 74554 96596 74556
rect 96620 74554 96676 74556
rect 96380 74502 96426 74554
rect 96426 74502 96436 74554
rect 96460 74502 96490 74554
rect 96490 74502 96502 74554
rect 96502 74502 96516 74554
rect 96540 74502 96554 74554
rect 96554 74502 96566 74554
rect 96566 74502 96596 74554
rect 96620 74502 96630 74554
rect 96630 74502 96676 74554
rect 96380 74500 96436 74502
rect 96460 74500 96516 74502
rect 96540 74500 96596 74502
rect 96620 74500 96676 74502
rect 97040 74010 97096 74012
rect 97120 74010 97176 74012
rect 97200 74010 97256 74012
rect 97280 74010 97336 74012
rect 97040 73958 97086 74010
rect 97086 73958 97096 74010
rect 97120 73958 97150 74010
rect 97150 73958 97162 74010
rect 97162 73958 97176 74010
rect 97200 73958 97214 74010
rect 97214 73958 97226 74010
rect 97226 73958 97256 74010
rect 97280 73958 97290 74010
rect 97290 73958 97336 74010
rect 97040 73956 97096 73958
rect 97120 73956 97176 73958
rect 97200 73956 97256 73958
rect 97280 73956 97336 73958
rect 96380 73466 96436 73468
rect 96460 73466 96516 73468
rect 96540 73466 96596 73468
rect 96620 73466 96676 73468
rect 96380 73414 96426 73466
rect 96426 73414 96436 73466
rect 96460 73414 96490 73466
rect 96490 73414 96502 73466
rect 96502 73414 96516 73466
rect 96540 73414 96554 73466
rect 96554 73414 96566 73466
rect 96566 73414 96596 73466
rect 96620 73414 96630 73466
rect 96630 73414 96676 73466
rect 96380 73412 96436 73414
rect 96460 73412 96516 73414
rect 96540 73412 96596 73414
rect 96620 73412 96676 73414
rect 97040 72922 97096 72924
rect 97120 72922 97176 72924
rect 97200 72922 97256 72924
rect 97280 72922 97336 72924
rect 97040 72870 97086 72922
rect 97086 72870 97096 72922
rect 97120 72870 97150 72922
rect 97150 72870 97162 72922
rect 97162 72870 97176 72922
rect 97200 72870 97214 72922
rect 97214 72870 97226 72922
rect 97226 72870 97256 72922
rect 97280 72870 97290 72922
rect 97290 72870 97336 72922
rect 97040 72868 97096 72870
rect 97120 72868 97176 72870
rect 97200 72868 97256 72870
rect 97280 72868 97336 72870
rect 96380 72378 96436 72380
rect 96460 72378 96516 72380
rect 96540 72378 96596 72380
rect 96620 72378 96676 72380
rect 96380 72326 96426 72378
rect 96426 72326 96436 72378
rect 96460 72326 96490 72378
rect 96490 72326 96502 72378
rect 96502 72326 96516 72378
rect 96540 72326 96554 72378
rect 96554 72326 96566 72378
rect 96566 72326 96596 72378
rect 96620 72326 96630 72378
rect 96630 72326 96676 72378
rect 96380 72324 96436 72326
rect 96460 72324 96516 72326
rect 96540 72324 96596 72326
rect 96620 72324 96676 72326
rect 97040 71834 97096 71836
rect 97120 71834 97176 71836
rect 97200 71834 97256 71836
rect 97280 71834 97336 71836
rect 97040 71782 97086 71834
rect 97086 71782 97096 71834
rect 97120 71782 97150 71834
rect 97150 71782 97162 71834
rect 97162 71782 97176 71834
rect 97200 71782 97214 71834
rect 97214 71782 97226 71834
rect 97226 71782 97256 71834
rect 97280 71782 97290 71834
rect 97290 71782 97336 71834
rect 97040 71780 97096 71782
rect 97120 71780 97176 71782
rect 97200 71780 97256 71782
rect 97280 71780 97336 71782
rect 96380 71290 96436 71292
rect 96460 71290 96516 71292
rect 96540 71290 96596 71292
rect 96620 71290 96676 71292
rect 96380 71238 96426 71290
rect 96426 71238 96436 71290
rect 96460 71238 96490 71290
rect 96490 71238 96502 71290
rect 96502 71238 96516 71290
rect 96540 71238 96554 71290
rect 96554 71238 96566 71290
rect 96566 71238 96596 71290
rect 96620 71238 96630 71290
rect 96630 71238 96676 71290
rect 96380 71236 96436 71238
rect 96460 71236 96516 71238
rect 96540 71236 96596 71238
rect 96620 71236 96676 71238
rect 97040 70746 97096 70748
rect 97120 70746 97176 70748
rect 97200 70746 97256 70748
rect 97280 70746 97336 70748
rect 97040 70694 97086 70746
rect 97086 70694 97096 70746
rect 97120 70694 97150 70746
rect 97150 70694 97162 70746
rect 97162 70694 97176 70746
rect 97200 70694 97214 70746
rect 97214 70694 97226 70746
rect 97226 70694 97256 70746
rect 97280 70694 97290 70746
rect 97290 70694 97336 70746
rect 97040 70692 97096 70694
rect 97120 70692 97176 70694
rect 97200 70692 97256 70694
rect 97280 70692 97336 70694
rect 96380 70202 96436 70204
rect 96460 70202 96516 70204
rect 96540 70202 96596 70204
rect 96620 70202 96676 70204
rect 96380 70150 96426 70202
rect 96426 70150 96436 70202
rect 96460 70150 96490 70202
rect 96490 70150 96502 70202
rect 96502 70150 96516 70202
rect 96540 70150 96554 70202
rect 96554 70150 96566 70202
rect 96566 70150 96596 70202
rect 96620 70150 96630 70202
rect 96630 70150 96676 70202
rect 96380 70148 96436 70150
rect 96460 70148 96516 70150
rect 96540 70148 96596 70150
rect 96620 70148 96676 70150
rect 97040 69658 97096 69660
rect 97120 69658 97176 69660
rect 97200 69658 97256 69660
rect 97280 69658 97336 69660
rect 97040 69606 97086 69658
rect 97086 69606 97096 69658
rect 97120 69606 97150 69658
rect 97150 69606 97162 69658
rect 97162 69606 97176 69658
rect 97200 69606 97214 69658
rect 97214 69606 97226 69658
rect 97226 69606 97256 69658
rect 97280 69606 97290 69658
rect 97290 69606 97336 69658
rect 97040 69604 97096 69606
rect 97120 69604 97176 69606
rect 97200 69604 97256 69606
rect 97280 69604 97336 69606
rect 96380 69114 96436 69116
rect 96460 69114 96516 69116
rect 96540 69114 96596 69116
rect 96620 69114 96676 69116
rect 96380 69062 96426 69114
rect 96426 69062 96436 69114
rect 96460 69062 96490 69114
rect 96490 69062 96502 69114
rect 96502 69062 96516 69114
rect 96540 69062 96554 69114
rect 96554 69062 96566 69114
rect 96566 69062 96596 69114
rect 96620 69062 96630 69114
rect 96630 69062 96676 69114
rect 96380 69060 96436 69062
rect 96460 69060 96516 69062
rect 96540 69060 96596 69062
rect 96620 69060 96676 69062
rect 97040 68570 97096 68572
rect 97120 68570 97176 68572
rect 97200 68570 97256 68572
rect 97280 68570 97336 68572
rect 97040 68518 97086 68570
rect 97086 68518 97096 68570
rect 97120 68518 97150 68570
rect 97150 68518 97162 68570
rect 97162 68518 97176 68570
rect 97200 68518 97214 68570
rect 97214 68518 97226 68570
rect 97226 68518 97256 68570
rect 97280 68518 97290 68570
rect 97290 68518 97336 68570
rect 97040 68516 97096 68518
rect 97120 68516 97176 68518
rect 97200 68516 97256 68518
rect 97280 68516 97336 68518
rect 96380 68026 96436 68028
rect 96460 68026 96516 68028
rect 96540 68026 96596 68028
rect 96620 68026 96676 68028
rect 96380 67974 96426 68026
rect 96426 67974 96436 68026
rect 96460 67974 96490 68026
rect 96490 67974 96502 68026
rect 96502 67974 96516 68026
rect 96540 67974 96554 68026
rect 96554 67974 96566 68026
rect 96566 67974 96596 68026
rect 96620 67974 96630 68026
rect 96630 67974 96676 68026
rect 96380 67972 96436 67974
rect 96460 67972 96516 67974
rect 96540 67972 96596 67974
rect 96620 67972 96676 67974
rect 97040 67482 97096 67484
rect 97120 67482 97176 67484
rect 97200 67482 97256 67484
rect 97280 67482 97336 67484
rect 97040 67430 97086 67482
rect 97086 67430 97096 67482
rect 97120 67430 97150 67482
rect 97150 67430 97162 67482
rect 97162 67430 97176 67482
rect 97200 67430 97214 67482
rect 97214 67430 97226 67482
rect 97226 67430 97256 67482
rect 97280 67430 97290 67482
rect 97290 67430 97336 67482
rect 97040 67428 97096 67430
rect 97120 67428 97176 67430
rect 97200 67428 97256 67430
rect 97280 67428 97336 67430
rect 96380 66938 96436 66940
rect 96460 66938 96516 66940
rect 96540 66938 96596 66940
rect 96620 66938 96676 66940
rect 96380 66886 96426 66938
rect 96426 66886 96436 66938
rect 96460 66886 96490 66938
rect 96490 66886 96502 66938
rect 96502 66886 96516 66938
rect 96540 66886 96554 66938
rect 96554 66886 96566 66938
rect 96566 66886 96596 66938
rect 96620 66886 96630 66938
rect 96630 66886 96676 66938
rect 96380 66884 96436 66886
rect 96460 66884 96516 66886
rect 96540 66884 96596 66886
rect 96620 66884 96676 66886
rect 97040 66394 97096 66396
rect 97120 66394 97176 66396
rect 97200 66394 97256 66396
rect 97280 66394 97336 66396
rect 97040 66342 97086 66394
rect 97086 66342 97096 66394
rect 97120 66342 97150 66394
rect 97150 66342 97162 66394
rect 97162 66342 97176 66394
rect 97200 66342 97214 66394
rect 97214 66342 97226 66394
rect 97226 66342 97256 66394
rect 97280 66342 97290 66394
rect 97290 66342 97336 66394
rect 97040 66340 97096 66342
rect 97120 66340 97176 66342
rect 97200 66340 97256 66342
rect 97280 66340 97336 66342
rect 96380 65850 96436 65852
rect 96460 65850 96516 65852
rect 96540 65850 96596 65852
rect 96620 65850 96676 65852
rect 96380 65798 96426 65850
rect 96426 65798 96436 65850
rect 96460 65798 96490 65850
rect 96490 65798 96502 65850
rect 96502 65798 96516 65850
rect 96540 65798 96554 65850
rect 96554 65798 96566 65850
rect 96566 65798 96596 65850
rect 96620 65798 96630 65850
rect 96630 65798 96676 65850
rect 96380 65796 96436 65798
rect 96460 65796 96516 65798
rect 96540 65796 96596 65798
rect 96620 65796 96676 65798
rect 97040 65306 97096 65308
rect 97120 65306 97176 65308
rect 97200 65306 97256 65308
rect 97280 65306 97336 65308
rect 97040 65254 97086 65306
rect 97086 65254 97096 65306
rect 97120 65254 97150 65306
rect 97150 65254 97162 65306
rect 97162 65254 97176 65306
rect 97200 65254 97214 65306
rect 97214 65254 97226 65306
rect 97226 65254 97256 65306
rect 97280 65254 97290 65306
rect 97290 65254 97336 65306
rect 97040 65252 97096 65254
rect 97120 65252 97176 65254
rect 97200 65252 97256 65254
rect 97280 65252 97336 65254
rect 96380 64762 96436 64764
rect 96460 64762 96516 64764
rect 96540 64762 96596 64764
rect 96620 64762 96676 64764
rect 96380 64710 96426 64762
rect 96426 64710 96436 64762
rect 96460 64710 96490 64762
rect 96490 64710 96502 64762
rect 96502 64710 96516 64762
rect 96540 64710 96554 64762
rect 96554 64710 96566 64762
rect 96566 64710 96596 64762
rect 96620 64710 96630 64762
rect 96630 64710 96676 64762
rect 96380 64708 96436 64710
rect 96460 64708 96516 64710
rect 96540 64708 96596 64710
rect 96620 64708 96676 64710
rect 97040 64218 97096 64220
rect 97120 64218 97176 64220
rect 97200 64218 97256 64220
rect 97280 64218 97336 64220
rect 97040 64166 97086 64218
rect 97086 64166 97096 64218
rect 97120 64166 97150 64218
rect 97150 64166 97162 64218
rect 97162 64166 97176 64218
rect 97200 64166 97214 64218
rect 97214 64166 97226 64218
rect 97226 64166 97256 64218
rect 97280 64166 97290 64218
rect 97290 64166 97336 64218
rect 97040 64164 97096 64166
rect 97120 64164 97176 64166
rect 97200 64164 97256 64166
rect 97280 64164 97336 64166
rect 96380 63674 96436 63676
rect 96460 63674 96516 63676
rect 96540 63674 96596 63676
rect 96620 63674 96676 63676
rect 96380 63622 96426 63674
rect 96426 63622 96436 63674
rect 96460 63622 96490 63674
rect 96490 63622 96502 63674
rect 96502 63622 96516 63674
rect 96540 63622 96554 63674
rect 96554 63622 96566 63674
rect 96566 63622 96596 63674
rect 96620 63622 96630 63674
rect 96630 63622 96676 63674
rect 96380 63620 96436 63622
rect 96460 63620 96516 63622
rect 96540 63620 96596 63622
rect 96620 63620 96676 63622
rect 97040 63130 97096 63132
rect 97120 63130 97176 63132
rect 97200 63130 97256 63132
rect 97280 63130 97336 63132
rect 97040 63078 97086 63130
rect 97086 63078 97096 63130
rect 97120 63078 97150 63130
rect 97150 63078 97162 63130
rect 97162 63078 97176 63130
rect 97200 63078 97214 63130
rect 97214 63078 97226 63130
rect 97226 63078 97256 63130
rect 97280 63078 97290 63130
rect 97290 63078 97336 63130
rect 97040 63076 97096 63078
rect 97120 63076 97176 63078
rect 97200 63076 97256 63078
rect 97280 63076 97336 63078
rect 100390 62636 100392 62656
rect 100392 62636 100444 62656
rect 100444 62636 100446 62656
rect 100390 62600 100446 62636
rect 96380 62586 96436 62588
rect 96460 62586 96516 62588
rect 96540 62586 96596 62588
rect 96620 62586 96676 62588
rect 96380 62534 96426 62586
rect 96426 62534 96436 62586
rect 96460 62534 96490 62586
rect 96490 62534 96502 62586
rect 96502 62534 96516 62586
rect 96540 62534 96554 62586
rect 96554 62534 96566 62586
rect 96566 62534 96596 62586
rect 96620 62534 96630 62586
rect 96630 62534 96676 62586
rect 96380 62532 96436 62534
rect 96460 62532 96516 62534
rect 96540 62532 96596 62534
rect 96620 62532 96676 62534
rect 96380 61498 96436 61500
rect 96460 61498 96516 61500
rect 96540 61498 96596 61500
rect 96620 61498 96676 61500
rect 96380 61446 96426 61498
rect 96426 61446 96436 61498
rect 96460 61446 96490 61498
rect 96490 61446 96502 61498
rect 96502 61446 96516 61498
rect 96540 61446 96554 61498
rect 96554 61446 96566 61498
rect 96566 61446 96596 61498
rect 96620 61446 96630 61498
rect 96630 61446 96676 61498
rect 96380 61444 96436 61446
rect 96460 61444 96516 61446
rect 96540 61444 96596 61446
rect 96620 61444 96676 61446
rect 97040 62042 97096 62044
rect 97120 62042 97176 62044
rect 97200 62042 97256 62044
rect 97280 62042 97336 62044
rect 97040 61990 97086 62042
rect 97086 61990 97096 62042
rect 97120 61990 97150 62042
rect 97150 61990 97162 62042
rect 97162 61990 97176 62042
rect 97200 61990 97214 62042
rect 97214 61990 97226 62042
rect 97226 61990 97256 62042
rect 97280 61990 97290 62042
rect 97290 61990 97336 62042
rect 97040 61988 97096 61990
rect 97120 61988 97176 61990
rect 97200 61988 97256 61990
rect 97280 61988 97336 61990
rect 100390 61920 100446 61976
rect 79506 58656 79562 58712
rect 79138 58520 79194 58576
rect 29182 58112 29238 58168
rect 97040 60954 97096 60956
rect 97120 60954 97176 60956
rect 97200 60954 97256 60956
rect 97280 60954 97336 60956
rect 97040 60902 97086 60954
rect 97086 60902 97096 60954
rect 97120 60902 97150 60954
rect 97150 60902 97162 60954
rect 97162 60902 97176 60954
rect 97200 60902 97214 60954
rect 97214 60902 97226 60954
rect 97226 60902 97256 60954
rect 97280 60902 97290 60954
rect 97290 60902 97336 60954
rect 97040 60900 97096 60902
rect 97120 60900 97176 60902
rect 97200 60900 97256 60902
rect 97280 60900 97336 60902
rect 86130 58520 86186 58576
rect 86130 58112 86186 58168
rect 83922 57976 83978 58032
rect 96380 60410 96436 60412
rect 96460 60410 96516 60412
rect 96540 60410 96596 60412
rect 96620 60410 96676 60412
rect 96380 60358 96426 60410
rect 96426 60358 96436 60410
rect 96460 60358 96490 60410
rect 96490 60358 96502 60410
rect 96502 60358 96516 60410
rect 96540 60358 96554 60410
rect 96554 60358 96566 60410
rect 96566 60358 96596 60410
rect 96620 60358 96630 60410
rect 96630 60358 96676 60410
rect 96380 60356 96436 60358
rect 96460 60356 96516 60358
rect 96540 60356 96596 60358
rect 96620 60356 96676 60358
rect 98936 60410 98992 60412
rect 99016 60410 99072 60412
rect 99096 60410 99152 60412
rect 99176 60410 99232 60412
rect 98936 60358 98982 60410
rect 98982 60358 98992 60410
rect 99016 60358 99046 60410
rect 99046 60358 99058 60410
rect 99058 60358 99072 60410
rect 99096 60358 99110 60410
rect 99110 60358 99122 60410
rect 99122 60358 99152 60410
rect 99176 60358 99186 60410
rect 99186 60358 99232 60410
rect 98936 60356 98992 60358
rect 99016 60356 99072 60358
rect 99096 60356 99152 60358
rect 99176 60356 99232 60358
rect 100390 61240 100446 61296
rect 100390 60580 100446 60616
rect 100390 60560 100392 60580
rect 100392 60560 100444 60580
rect 100444 60560 100446 60580
rect 97040 59866 97096 59868
rect 97120 59866 97176 59868
rect 97200 59866 97256 59868
rect 97280 59866 97336 59868
rect 97040 59814 97086 59866
rect 97086 59814 97096 59866
rect 97120 59814 97150 59866
rect 97150 59814 97162 59866
rect 97162 59814 97176 59866
rect 97200 59814 97214 59866
rect 97214 59814 97226 59866
rect 97226 59814 97256 59866
rect 97280 59814 97290 59866
rect 97290 59814 97336 59866
rect 97040 59812 97096 59814
rect 97120 59812 97176 59814
rect 97200 59812 97256 59814
rect 97280 59812 97336 59814
rect 28170 57840 28226 57896
rect 81806 57840 81862 57896
rect 87878 57840 87934 57896
rect 97078 53760 97134 53816
rect 98274 58520 98330 58576
rect 100390 59916 100392 59936
rect 100392 59916 100444 59936
rect 100444 59916 100446 59936
rect 100390 59880 100446 59916
rect 99672 59866 99728 59868
rect 99752 59866 99808 59868
rect 99832 59866 99888 59868
rect 99912 59866 99968 59868
rect 99672 59814 99718 59866
rect 99718 59814 99728 59866
rect 99752 59814 99782 59866
rect 99782 59814 99794 59866
rect 99794 59814 99808 59866
rect 99832 59814 99846 59866
rect 99846 59814 99858 59866
rect 99858 59814 99888 59866
rect 99912 59814 99922 59866
rect 99922 59814 99968 59866
rect 99672 59812 99728 59814
rect 99752 59812 99808 59814
rect 99832 59812 99888 59814
rect 99912 59812 99968 59814
rect 98936 59322 98992 59324
rect 99016 59322 99072 59324
rect 99096 59322 99152 59324
rect 99176 59322 99232 59324
rect 98936 59270 98982 59322
rect 98982 59270 98992 59322
rect 99016 59270 99046 59322
rect 99046 59270 99058 59322
rect 99058 59270 99072 59322
rect 99096 59270 99110 59322
rect 99110 59270 99122 59322
rect 99122 59270 99152 59322
rect 99176 59270 99186 59322
rect 99186 59270 99232 59322
rect 98936 59268 98992 59270
rect 99016 59268 99072 59270
rect 99096 59268 99152 59270
rect 99176 59268 99232 59270
rect 99672 58778 99728 58780
rect 99752 58778 99808 58780
rect 99832 58778 99888 58780
rect 99912 58778 99968 58780
rect 99672 58726 99718 58778
rect 99718 58726 99728 58778
rect 99752 58726 99782 58778
rect 99782 58726 99794 58778
rect 99794 58726 99808 58778
rect 99832 58726 99846 58778
rect 99846 58726 99858 58778
rect 99858 58726 99888 58778
rect 99912 58726 99922 58778
rect 99922 58726 99968 58778
rect 99672 58724 99728 58726
rect 99752 58724 99808 58726
rect 99832 58724 99888 58726
rect 99912 58724 99968 58726
rect 98936 58234 98992 58236
rect 99016 58234 99072 58236
rect 99096 58234 99152 58236
rect 99176 58234 99232 58236
rect 98936 58182 98982 58234
rect 98982 58182 98992 58234
rect 99016 58182 99046 58234
rect 99046 58182 99058 58234
rect 99058 58182 99072 58234
rect 99096 58182 99110 58234
rect 99110 58182 99122 58234
rect 99122 58182 99152 58234
rect 99176 58182 99186 58234
rect 99186 58182 99232 58234
rect 98936 58180 98992 58182
rect 99016 58180 99072 58182
rect 99096 58180 99152 58182
rect 99176 58180 99232 58182
rect 100114 57840 100170 57896
rect 99672 57690 99728 57692
rect 99752 57690 99808 57692
rect 99832 57690 99888 57692
rect 99912 57690 99968 57692
rect 99672 57638 99718 57690
rect 99718 57638 99728 57690
rect 99752 57638 99782 57690
rect 99782 57638 99794 57690
rect 99794 57638 99808 57690
rect 99832 57638 99846 57690
rect 99846 57638 99858 57690
rect 99858 57638 99888 57690
rect 99912 57638 99922 57690
rect 99922 57638 99968 57690
rect 99672 57636 99728 57638
rect 99752 57636 99808 57638
rect 99832 57636 99888 57638
rect 99912 57636 99968 57638
rect 98936 57146 98992 57148
rect 99016 57146 99072 57148
rect 99096 57146 99152 57148
rect 99176 57146 99232 57148
rect 98936 57094 98982 57146
rect 98982 57094 98992 57146
rect 99016 57094 99046 57146
rect 99046 57094 99058 57146
rect 99058 57094 99072 57146
rect 99096 57094 99110 57146
rect 99110 57094 99122 57146
rect 99122 57094 99152 57146
rect 99176 57094 99186 57146
rect 99186 57094 99232 57146
rect 98936 57092 98992 57094
rect 99016 57092 99072 57094
rect 99096 57092 99152 57094
rect 99176 57092 99232 57094
rect 99672 56602 99728 56604
rect 99752 56602 99808 56604
rect 99832 56602 99888 56604
rect 99912 56602 99968 56604
rect 99672 56550 99718 56602
rect 99718 56550 99728 56602
rect 99752 56550 99782 56602
rect 99782 56550 99794 56602
rect 99794 56550 99808 56602
rect 99832 56550 99846 56602
rect 99846 56550 99858 56602
rect 99858 56550 99888 56602
rect 99912 56550 99922 56602
rect 99922 56550 99968 56602
rect 99672 56548 99728 56550
rect 99752 56548 99808 56550
rect 99832 56548 99888 56550
rect 99912 56548 99968 56550
rect 98936 56058 98992 56060
rect 99016 56058 99072 56060
rect 99096 56058 99152 56060
rect 99176 56058 99232 56060
rect 98936 56006 98982 56058
rect 98982 56006 98992 56058
rect 99016 56006 99046 56058
rect 99046 56006 99058 56058
rect 99058 56006 99072 56058
rect 99096 56006 99110 56058
rect 99110 56006 99122 56058
rect 99122 56006 99152 56058
rect 99176 56006 99186 56058
rect 99186 56006 99232 56058
rect 98936 56004 98992 56006
rect 99016 56004 99072 56006
rect 99096 56004 99152 56006
rect 99176 56004 99232 56006
rect 99672 55514 99728 55516
rect 99752 55514 99808 55516
rect 99832 55514 99888 55516
rect 99912 55514 99968 55516
rect 99672 55462 99718 55514
rect 99718 55462 99728 55514
rect 99752 55462 99782 55514
rect 99782 55462 99794 55514
rect 99794 55462 99808 55514
rect 99832 55462 99846 55514
rect 99846 55462 99858 55514
rect 99858 55462 99888 55514
rect 99912 55462 99922 55514
rect 99922 55462 99968 55514
rect 99672 55460 99728 55462
rect 99752 55460 99808 55462
rect 99832 55460 99888 55462
rect 99912 55460 99968 55462
rect 98936 54970 98992 54972
rect 99016 54970 99072 54972
rect 99096 54970 99152 54972
rect 99176 54970 99232 54972
rect 98936 54918 98982 54970
rect 98982 54918 98992 54970
rect 99016 54918 99046 54970
rect 99046 54918 99058 54970
rect 99058 54918 99072 54970
rect 99096 54918 99110 54970
rect 99110 54918 99122 54970
rect 99122 54918 99152 54970
rect 99176 54918 99186 54970
rect 99186 54918 99232 54970
rect 98936 54916 98992 54918
rect 99016 54916 99072 54918
rect 99096 54916 99152 54918
rect 99176 54916 99232 54918
rect 99672 54426 99728 54428
rect 99752 54426 99808 54428
rect 99832 54426 99888 54428
rect 99912 54426 99968 54428
rect 99672 54374 99718 54426
rect 99718 54374 99728 54426
rect 99752 54374 99782 54426
rect 99782 54374 99794 54426
rect 99794 54374 99808 54426
rect 99832 54374 99846 54426
rect 99846 54374 99858 54426
rect 99858 54374 99888 54426
rect 99912 54374 99922 54426
rect 99922 54374 99968 54426
rect 99672 54372 99728 54374
rect 99752 54372 99808 54374
rect 99832 54372 99888 54374
rect 99912 54372 99968 54374
rect 98936 53882 98992 53884
rect 99016 53882 99072 53884
rect 99096 53882 99152 53884
rect 99176 53882 99232 53884
rect 98936 53830 98982 53882
rect 98982 53830 98992 53882
rect 99016 53830 99046 53882
rect 99046 53830 99058 53882
rect 99058 53830 99072 53882
rect 99096 53830 99110 53882
rect 99110 53830 99122 53882
rect 99122 53830 99152 53882
rect 99176 53830 99186 53882
rect 99186 53830 99232 53882
rect 98936 53828 98992 53830
rect 99016 53828 99072 53830
rect 99096 53828 99152 53830
rect 99176 53828 99232 53830
rect 99672 53338 99728 53340
rect 99752 53338 99808 53340
rect 99832 53338 99888 53340
rect 99912 53338 99968 53340
rect 99672 53286 99718 53338
rect 99718 53286 99728 53338
rect 99752 53286 99782 53338
rect 99782 53286 99794 53338
rect 99794 53286 99808 53338
rect 99832 53286 99846 53338
rect 99846 53286 99858 53338
rect 99858 53286 99888 53338
rect 99912 53286 99922 53338
rect 99922 53286 99968 53338
rect 99672 53284 99728 53286
rect 99752 53284 99808 53286
rect 99832 53284 99888 53286
rect 99912 53284 99968 53286
rect 98936 52794 98992 52796
rect 99016 52794 99072 52796
rect 99096 52794 99152 52796
rect 99176 52794 99232 52796
rect 98936 52742 98982 52794
rect 98982 52742 98992 52794
rect 99016 52742 99046 52794
rect 99046 52742 99058 52794
rect 99058 52742 99072 52794
rect 99096 52742 99110 52794
rect 99110 52742 99122 52794
rect 99122 52742 99152 52794
rect 99176 52742 99186 52794
rect 99186 52742 99232 52794
rect 98936 52740 98992 52742
rect 99016 52740 99072 52742
rect 99096 52740 99152 52742
rect 99176 52740 99232 52742
rect 99672 52250 99728 52252
rect 99752 52250 99808 52252
rect 99832 52250 99888 52252
rect 99912 52250 99968 52252
rect 99672 52198 99718 52250
rect 99718 52198 99728 52250
rect 99752 52198 99782 52250
rect 99782 52198 99794 52250
rect 99794 52198 99808 52250
rect 99832 52198 99846 52250
rect 99846 52198 99858 52250
rect 99858 52198 99888 52250
rect 99912 52198 99922 52250
rect 99922 52198 99968 52250
rect 99672 52196 99728 52198
rect 99752 52196 99808 52198
rect 99832 52196 99888 52198
rect 99912 52196 99968 52198
rect 98936 51706 98992 51708
rect 99016 51706 99072 51708
rect 99096 51706 99152 51708
rect 99176 51706 99232 51708
rect 98936 51654 98982 51706
rect 98982 51654 98992 51706
rect 99016 51654 99046 51706
rect 99046 51654 99058 51706
rect 99058 51654 99072 51706
rect 99096 51654 99110 51706
rect 99110 51654 99122 51706
rect 99122 51654 99152 51706
rect 99176 51654 99186 51706
rect 99186 51654 99232 51706
rect 98936 51652 98992 51654
rect 99016 51652 99072 51654
rect 99096 51652 99152 51654
rect 99176 51652 99232 51654
rect 99672 51162 99728 51164
rect 99752 51162 99808 51164
rect 99832 51162 99888 51164
rect 99912 51162 99968 51164
rect 99672 51110 99718 51162
rect 99718 51110 99728 51162
rect 99752 51110 99782 51162
rect 99782 51110 99794 51162
rect 99794 51110 99808 51162
rect 99832 51110 99846 51162
rect 99846 51110 99858 51162
rect 99858 51110 99888 51162
rect 99912 51110 99922 51162
rect 99922 51110 99968 51162
rect 99672 51108 99728 51110
rect 99752 51108 99808 51110
rect 99832 51108 99888 51110
rect 99912 51108 99968 51110
rect 98936 50618 98992 50620
rect 99016 50618 99072 50620
rect 99096 50618 99152 50620
rect 99176 50618 99232 50620
rect 98936 50566 98982 50618
rect 98982 50566 98992 50618
rect 99016 50566 99046 50618
rect 99046 50566 99058 50618
rect 99058 50566 99072 50618
rect 99096 50566 99110 50618
rect 99110 50566 99122 50618
rect 99122 50566 99152 50618
rect 99176 50566 99186 50618
rect 99186 50566 99232 50618
rect 98936 50564 98992 50566
rect 99016 50564 99072 50566
rect 99096 50564 99152 50566
rect 99176 50564 99232 50566
rect 99672 50074 99728 50076
rect 99752 50074 99808 50076
rect 99832 50074 99888 50076
rect 99912 50074 99968 50076
rect 99672 50022 99718 50074
rect 99718 50022 99728 50074
rect 99752 50022 99782 50074
rect 99782 50022 99794 50074
rect 99794 50022 99808 50074
rect 99832 50022 99846 50074
rect 99846 50022 99858 50074
rect 99858 50022 99888 50074
rect 99912 50022 99922 50074
rect 99922 50022 99968 50074
rect 99672 50020 99728 50022
rect 99752 50020 99808 50022
rect 99832 50020 99888 50022
rect 99912 50020 99968 50022
rect 98936 49530 98992 49532
rect 99016 49530 99072 49532
rect 99096 49530 99152 49532
rect 99176 49530 99232 49532
rect 98936 49478 98982 49530
rect 98982 49478 98992 49530
rect 99016 49478 99046 49530
rect 99046 49478 99058 49530
rect 99058 49478 99072 49530
rect 99096 49478 99110 49530
rect 99110 49478 99122 49530
rect 99122 49478 99152 49530
rect 99176 49478 99186 49530
rect 99186 49478 99232 49530
rect 98936 49476 98992 49478
rect 99016 49476 99072 49478
rect 99096 49476 99152 49478
rect 99176 49476 99232 49478
rect 99672 48986 99728 48988
rect 99752 48986 99808 48988
rect 99832 48986 99888 48988
rect 99912 48986 99968 48988
rect 99672 48934 99718 48986
rect 99718 48934 99728 48986
rect 99752 48934 99782 48986
rect 99782 48934 99794 48986
rect 99794 48934 99808 48986
rect 99832 48934 99846 48986
rect 99846 48934 99858 48986
rect 99858 48934 99888 48986
rect 99912 48934 99922 48986
rect 99922 48934 99968 48986
rect 99672 48932 99728 48934
rect 99752 48932 99808 48934
rect 99832 48932 99888 48934
rect 99912 48932 99968 48934
rect 98936 48442 98992 48444
rect 99016 48442 99072 48444
rect 99096 48442 99152 48444
rect 99176 48442 99232 48444
rect 98936 48390 98982 48442
rect 98982 48390 98992 48442
rect 99016 48390 99046 48442
rect 99046 48390 99058 48442
rect 99058 48390 99072 48442
rect 99096 48390 99110 48442
rect 99110 48390 99122 48442
rect 99122 48390 99152 48442
rect 99176 48390 99186 48442
rect 99186 48390 99232 48442
rect 98936 48388 98992 48390
rect 99016 48388 99072 48390
rect 99096 48388 99152 48390
rect 99176 48388 99232 48390
rect 99672 47898 99728 47900
rect 99752 47898 99808 47900
rect 99832 47898 99888 47900
rect 99912 47898 99968 47900
rect 99672 47846 99718 47898
rect 99718 47846 99728 47898
rect 99752 47846 99782 47898
rect 99782 47846 99794 47898
rect 99794 47846 99808 47898
rect 99832 47846 99846 47898
rect 99846 47846 99858 47898
rect 99858 47846 99888 47898
rect 99912 47846 99922 47898
rect 99922 47846 99968 47898
rect 99672 47844 99728 47846
rect 99752 47844 99808 47846
rect 99832 47844 99888 47846
rect 99912 47844 99968 47846
rect 98936 47354 98992 47356
rect 99016 47354 99072 47356
rect 99096 47354 99152 47356
rect 99176 47354 99232 47356
rect 98936 47302 98982 47354
rect 98982 47302 98992 47354
rect 99016 47302 99046 47354
rect 99046 47302 99058 47354
rect 99058 47302 99072 47354
rect 99096 47302 99110 47354
rect 99110 47302 99122 47354
rect 99122 47302 99152 47354
rect 99176 47302 99186 47354
rect 99186 47302 99232 47354
rect 98936 47300 98992 47302
rect 99016 47300 99072 47302
rect 99096 47300 99152 47302
rect 99176 47300 99232 47302
rect 99672 46810 99728 46812
rect 99752 46810 99808 46812
rect 99832 46810 99888 46812
rect 99912 46810 99968 46812
rect 99672 46758 99718 46810
rect 99718 46758 99728 46810
rect 99752 46758 99782 46810
rect 99782 46758 99794 46810
rect 99794 46758 99808 46810
rect 99832 46758 99846 46810
rect 99846 46758 99858 46810
rect 99858 46758 99888 46810
rect 99912 46758 99922 46810
rect 99922 46758 99968 46810
rect 99672 46756 99728 46758
rect 99752 46756 99808 46758
rect 99832 46756 99888 46758
rect 99912 46756 99968 46758
rect 98936 46266 98992 46268
rect 99016 46266 99072 46268
rect 99096 46266 99152 46268
rect 99176 46266 99232 46268
rect 98936 46214 98982 46266
rect 98982 46214 98992 46266
rect 99016 46214 99046 46266
rect 99046 46214 99058 46266
rect 99058 46214 99072 46266
rect 99096 46214 99110 46266
rect 99110 46214 99122 46266
rect 99122 46214 99152 46266
rect 99176 46214 99186 46266
rect 99186 46214 99232 46266
rect 98936 46212 98992 46214
rect 99016 46212 99072 46214
rect 99096 46212 99152 46214
rect 99176 46212 99232 46214
rect 97262 4120 97318 4176
rect 2686 3848 2742 3904
rect 1312 3834 1368 3836
rect 1392 3834 1448 3836
rect 1312 3782 1322 3834
rect 1322 3782 1368 3834
rect 1392 3782 1438 3834
rect 1438 3782 1448 3834
rect 1312 3780 1368 3782
rect 1392 3780 1448 3782
rect 99672 45722 99728 45724
rect 99752 45722 99808 45724
rect 99832 45722 99888 45724
rect 99912 45722 99968 45724
rect 99672 45670 99718 45722
rect 99718 45670 99728 45722
rect 99752 45670 99782 45722
rect 99782 45670 99794 45722
rect 99794 45670 99808 45722
rect 99832 45670 99846 45722
rect 99846 45670 99858 45722
rect 99858 45670 99888 45722
rect 99912 45670 99922 45722
rect 99922 45670 99968 45722
rect 99672 45668 99728 45670
rect 99752 45668 99808 45670
rect 99832 45668 99888 45670
rect 99912 45668 99968 45670
rect 98936 45178 98992 45180
rect 99016 45178 99072 45180
rect 99096 45178 99152 45180
rect 99176 45178 99232 45180
rect 98936 45126 98982 45178
rect 98982 45126 98992 45178
rect 99016 45126 99046 45178
rect 99046 45126 99058 45178
rect 99058 45126 99072 45178
rect 99096 45126 99110 45178
rect 99110 45126 99122 45178
rect 99122 45126 99152 45178
rect 99176 45126 99186 45178
rect 99186 45126 99232 45178
rect 98936 45124 98992 45126
rect 99016 45124 99072 45126
rect 99096 45124 99152 45126
rect 99176 45124 99232 45126
rect 99672 44634 99728 44636
rect 99752 44634 99808 44636
rect 99832 44634 99888 44636
rect 99912 44634 99968 44636
rect 99672 44582 99718 44634
rect 99718 44582 99728 44634
rect 99752 44582 99782 44634
rect 99782 44582 99794 44634
rect 99794 44582 99808 44634
rect 99832 44582 99846 44634
rect 99846 44582 99858 44634
rect 99858 44582 99888 44634
rect 99912 44582 99922 44634
rect 99922 44582 99968 44634
rect 99672 44580 99728 44582
rect 99752 44580 99808 44582
rect 99832 44580 99888 44582
rect 99912 44580 99968 44582
rect 98936 44090 98992 44092
rect 99016 44090 99072 44092
rect 99096 44090 99152 44092
rect 99176 44090 99232 44092
rect 98936 44038 98982 44090
rect 98982 44038 98992 44090
rect 99016 44038 99046 44090
rect 99046 44038 99058 44090
rect 99058 44038 99072 44090
rect 99096 44038 99110 44090
rect 99110 44038 99122 44090
rect 99122 44038 99152 44090
rect 99176 44038 99186 44090
rect 99186 44038 99232 44090
rect 98936 44036 98992 44038
rect 99016 44036 99072 44038
rect 99096 44036 99152 44038
rect 99176 44036 99232 44038
rect 99672 43546 99728 43548
rect 99752 43546 99808 43548
rect 99832 43546 99888 43548
rect 99912 43546 99968 43548
rect 99672 43494 99718 43546
rect 99718 43494 99728 43546
rect 99752 43494 99782 43546
rect 99782 43494 99794 43546
rect 99794 43494 99808 43546
rect 99832 43494 99846 43546
rect 99846 43494 99858 43546
rect 99858 43494 99888 43546
rect 99912 43494 99922 43546
rect 99922 43494 99968 43546
rect 99672 43492 99728 43494
rect 99752 43492 99808 43494
rect 99832 43492 99888 43494
rect 99912 43492 99968 43494
rect 98936 43002 98992 43004
rect 99016 43002 99072 43004
rect 99096 43002 99152 43004
rect 99176 43002 99232 43004
rect 98936 42950 98982 43002
rect 98982 42950 98992 43002
rect 99016 42950 99046 43002
rect 99046 42950 99058 43002
rect 99058 42950 99072 43002
rect 99096 42950 99110 43002
rect 99110 42950 99122 43002
rect 99122 42950 99152 43002
rect 99176 42950 99186 43002
rect 99186 42950 99232 43002
rect 98936 42948 98992 42950
rect 99016 42948 99072 42950
rect 99096 42948 99152 42950
rect 99176 42948 99232 42950
rect 99672 42458 99728 42460
rect 99752 42458 99808 42460
rect 99832 42458 99888 42460
rect 99912 42458 99968 42460
rect 99672 42406 99718 42458
rect 99718 42406 99728 42458
rect 99752 42406 99782 42458
rect 99782 42406 99794 42458
rect 99794 42406 99808 42458
rect 99832 42406 99846 42458
rect 99846 42406 99858 42458
rect 99858 42406 99888 42458
rect 99912 42406 99922 42458
rect 99922 42406 99968 42458
rect 99672 42404 99728 42406
rect 99752 42404 99808 42406
rect 99832 42404 99888 42406
rect 99912 42404 99968 42406
rect 98936 41914 98992 41916
rect 99016 41914 99072 41916
rect 99096 41914 99152 41916
rect 99176 41914 99232 41916
rect 98936 41862 98982 41914
rect 98982 41862 98992 41914
rect 99016 41862 99046 41914
rect 99046 41862 99058 41914
rect 99058 41862 99072 41914
rect 99096 41862 99110 41914
rect 99110 41862 99122 41914
rect 99122 41862 99152 41914
rect 99176 41862 99186 41914
rect 99186 41862 99232 41914
rect 98936 41860 98992 41862
rect 99016 41860 99072 41862
rect 99096 41860 99152 41862
rect 99176 41860 99232 41862
rect 99672 41370 99728 41372
rect 99752 41370 99808 41372
rect 99832 41370 99888 41372
rect 99912 41370 99968 41372
rect 99672 41318 99718 41370
rect 99718 41318 99728 41370
rect 99752 41318 99782 41370
rect 99782 41318 99794 41370
rect 99794 41318 99808 41370
rect 99832 41318 99846 41370
rect 99846 41318 99858 41370
rect 99858 41318 99888 41370
rect 99912 41318 99922 41370
rect 99922 41318 99968 41370
rect 99672 41316 99728 41318
rect 99752 41316 99808 41318
rect 99832 41316 99888 41318
rect 99912 41316 99968 41318
rect 98936 40826 98992 40828
rect 99016 40826 99072 40828
rect 99096 40826 99152 40828
rect 99176 40826 99232 40828
rect 98936 40774 98982 40826
rect 98982 40774 98992 40826
rect 99016 40774 99046 40826
rect 99046 40774 99058 40826
rect 99058 40774 99072 40826
rect 99096 40774 99110 40826
rect 99110 40774 99122 40826
rect 99122 40774 99152 40826
rect 99176 40774 99186 40826
rect 99186 40774 99232 40826
rect 98936 40772 98992 40774
rect 99016 40772 99072 40774
rect 99096 40772 99152 40774
rect 99176 40772 99232 40774
rect 99672 40282 99728 40284
rect 99752 40282 99808 40284
rect 99832 40282 99888 40284
rect 99912 40282 99968 40284
rect 99672 40230 99718 40282
rect 99718 40230 99728 40282
rect 99752 40230 99782 40282
rect 99782 40230 99794 40282
rect 99794 40230 99808 40282
rect 99832 40230 99846 40282
rect 99846 40230 99858 40282
rect 99858 40230 99888 40282
rect 99912 40230 99922 40282
rect 99922 40230 99968 40282
rect 99672 40228 99728 40230
rect 99752 40228 99808 40230
rect 99832 40228 99888 40230
rect 99912 40228 99968 40230
rect 98936 39738 98992 39740
rect 99016 39738 99072 39740
rect 99096 39738 99152 39740
rect 99176 39738 99232 39740
rect 98936 39686 98982 39738
rect 98982 39686 98992 39738
rect 99016 39686 99046 39738
rect 99046 39686 99058 39738
rect 99058 39686 99072 39738
rect 99096 39686 99110 39738
rect 99110 39686 99122 39738
rect 99122 39686 99152 39738
rect 99176 39686 99186 39738
rect 99186 39686 99232 39738
rect 98936 39684 98992 39686
rect 99016 39684 99072 39686
rect 99096 39684 99152 39686
rect 99176 39684 99232 39686
rect 99672 39194 99728 39196
rect 99752 39194 99808 39196
rect 99832 39194 99888 39196
rect 99912 39194 99968 39196
rect 99672 39142 99718 39194
rect 99718 39142 99728 39194
rect 99752 39142 99782 39194
rect 99782 39142 99794 39194
rect 99794 39142 99808 39194
rect 99832 39142 99846 39194
rect 99846 39142 99858 39194
rect 99858 39142 99888 39194
rect 99912 39142 99922 39194
rect 99922 39142 99968 39194
rect 99672 39140 99728 39142
rect 99752 39140 99808 39142
rect 99832 39140 99888 39142
rect 99912 39140 99968 39142
rect 98936 38650 98992 38652
rect 99016 38650 99072 38652
rect 99096 38650 99152 38652
rect 99176 38650 99232 38652
rect 98936 38598 98982 38650
rect 98982 38598 98992 38650
rect 99016 38598 99046 38650
rect 99046 38598 99058 38650
rect 99058 38598 99072 38650
rect 99096 38598 99110 38650
rect 99110 38598 99122 38650
rect 99122 38598 99152 38650
rect 99176 38598 99186 38650
rect 99186 38598 99232 38650
rect 98936 38596 98992 38598
rect 99016 38596 99072 38598
rect 99096 38596 99152 38598
rect 99176 38596 99232 38598
rect 99672 38106 99728 38108
rect 99752 38106 99808 38108
rect 99832 38106 99888 38108
rect 99912 38106 99968 38108
rect 99672 38054 99718 38106
rect 99718 38054 99728 38106
rect 99752 38054 99782 38106
rect 99782 38054 99794 38106
rect 99794 38054 99808 38106
rect 99832 38054 99846 38106
rect 99846 38054 99858 38106
rect 99858 38054 99888 38106
rect 99912 38054 99922 38106
rect 99922 38054 99968 38106
rect 99672 38052 99728 38054
rect 99752 38052 99808 38054
rect 99832 38052 99888 38054
rect 99912 38052 99968 38054
rect 98936 37562 98992 37564
rect 99016 37562 99072 37564
rect 99096 37562 99152 37564
rect 99176 37562 99232 37564
rect 98936 37510 98982 37562
rect 98982 37510 98992 37562
rect 99016 37510 99046 37562
rect 99046 37510 99058 37562
rect 99058 37510 99072 37562
rect 99096 37510 99110 37562
rect 99110 37510 99122 37562
rect 99122 37510 99152 37562
rect 99176 37510 99186 37562
rect 99186 37510 99232 37562
rect 98936 37508 98992 37510
rect 99016 37508 99072 37510
rect 99096 37508 99152 37510
rect 99176 37508 99232 37510
rect 99672 37018 99728 37020
rect 99752 37018 99808 37020
rect 99832 37018 99888 37020
rect 99912 37018 99968 37020
rect 99672 36966 99718 37018
rect 99718 36966 99728 37018
rect 99752 36966 99782 37018
rect 99782 36966 99794 37018
rect 99794 36966 99808 37018
rect 99832 36966 99846 37018
rect 99846 36966 99858 37018
rect 99858 36966 99888 37018
rect 99912 36966 99922 37018
rect 99922 36966 99968 37018
rect 99672 36964 99728 36966
rect 99752 36964 99808 36966
rect 99832 36964 99888 36966
rect 99912 36964 99968 36966
rect 98936 36474 98992 36476
rect 99016 36474 99072 36476
rect 99096 36474 99152 36476
rect 99176 36474 99232 36476
rect 98936 36422 98982 36474
rect 98982 36422 98992 36474
rect 99016 36422 99046 36474
rect 99046 36422 99058 36474
rect 99058 36422 99072 36474
rect 99096 36422 99110 36474
rect 99110 36422 99122 36474
rect 99122 36422 99152 36474
rect 99176 36422 99186 36474
rect 99186 36422 99232 36474
rect 98936 36420 98992 36422
rect 99016 36420 99072 36422
rect 99096 36420 99152 36422
rect 99176 36420 99232 36422
rect 99672 35930 99728 35932
rect 99752 35930 99808 35932
rect 99832 35930 99888 35932
rect 99912 35930 99968 35932
rect 99672 35878 99718 35930
rect 99718 35878 99728 35930
rect 99752 35878 99782 35930
rect 99782 35878 99794 35930
rect 99794 35878 99808 35930
rect 99832 35878 99846 35930
rect 99846 35878 99858 35930
rect 99858 35878 99888 35930
rect 99912 35878 99922 35930
rect 99922 35878 99968 35930
rect 99672 35876 99728 35878
rect 99752 35876 99808 35878
rect 99832 35876 99888 35878
rect 99912 35876 99968 35878
rect 98936 35386 98992 35388
rect 99016 35386 99072 35388
rect 99096 35386 99152 35388
rect 99176 35386 99232 35388
rect 98936 35334 98982 35386
rect 98982 35334 98992 35386
rect 99016 35334 99046 35386
rect 99046 35334 99058 35386
rect 99058 35334 99072 35386
rect 99096 35334 99110 35386
rect 99110 35334 99122 35386
rect 99122 35334 99152 35386
rect 99176 35334 99186 35386
rect 99186 35334 99232 35386
rect 98936 35332 98992 35334
rect 99016 35332 99072 35334
rect 99096 35332 99152 35334
rect 99176 35332 99232 35334
rect 99672 34842 99728 34844
rect 99752 34842 99808 34844
rect 99832 34842 99888 34844
rect 99912 34842 99968 34844
rect 99672 34790 99718 34842
rect 99718 34790 99728 34842
rect 99752 34790 99782 34842
rect 99782 34790 99794 34842
rect 99794 34790 99808 34842
rect 99832 34790 99846 34842
rect 99846 34790 99858 34842
rect 99858 34790 99888 34842
rect 99912 34790 99922 34842
rect 99922 34790 99968 34842
rect 99672 34788 99728 34790
rect 99752 34788 99808 34790
rect 99832 34788 99888 34790
rect 99912 34788 99968 34790
rect 98936 34298 98992 34300
rect 99016 34298 99072 34300
rect 99096 34298 99152 34300
rect 99176 34298 99232 34300
rect 98936 34246 98982 34298
rect 98982 34246 98992 34298
rect 99016 34246 99046 34298
rect 99046 34246 99058 34298
rect 99058 34246 99072 34298
rect 99096 34246 99110 34298
rect 99110 34246 99122 34298
rect 99122 34246 99152 34298
rect 99176 34246 99186 34298
rect 99186 34246 99232 34298
rect 98936 34244 98992 34246
rect 99016 34244 99072 34246
rect 99096 34244 99152 34246
rect 99176 34244 99232 34246
rect 99672 33754 99728 33756
rect 99752 33754 99808 33756
rect 99832 33754 99888 33756
rect 99912 33754 99968 33756
rect 99672 33702 99718 33754
rect 99718 33702 99728 33754
rect 99752 33702 99782 33754
rect 99782 33702 99794 33754
rect 99794 33702 99808 33754
rect 99832 33702 99846 33754
rect 99846 33702 99858 33754
rect 99858 33702 99888 33754
rect 99912 33702 99922 33754
rect 99922 33702 99968 33754
rect 99672 33700 99728 33702
rect 99752 33700 99808 33702
rect 99832 33700 99888 33702
rect 99912 33700 99968 33702
rect 98936 33210 98992 33212
rect 99016 33210 99072 33212
rect 99096 33210 99152 33212
rect 99176 33210 99232 33212
rect 98936 33158 98982 33210
rect 98982 33158 98992 33210
rect 99016 33158 99046 33210
rect 99046 33158 99058 33210
rect 99058 33158 99072 33210
rect 99096 33158 99110 33210
rect 99110 33158 99122 33210
rect 99122 33158 99152 33210
rect 99176 33158 99186 33210
rect 99186 33158 99232 33210
rect 98936 33156 98992 33158
rect 99016 33156 99072 33158
rect 99096 33156 99152 33158
rect 99176 33156 99232 33158
rect 99672 32666 99728 32668
rect 99752 32666 99808 32668
rect 99832 32666 99888 32668
rect 99912 32666 99968 32668
rect 99672 32614 99718 32666
rect 99718 32614 99728 32666
rect 99752 32614 99782 32666
rect 99782 32614 99794 32666
rect 99794 32614 99808 32666
rect 99832 32614 99846 32666
rect 99846 32614 99858 32666
rect 99858 32614 99888 32666
rect 99912 32614 99922 32666
rect 99922 32614 99968 32666
rect 99672 32612 99728 32614
rect 99752 32612 99808 32614
rect 99832 32612 99888 32614
rect 99912 32612 99968 32614
rect 98936 32122 98992 32124
rect 99016 32122 99072 32124
rect 99096 32122 99152 32124
rect 99176 32122 99232 32124
rect 98936 32070 98982 32122
rect 98982 32070 98992 32122
rect 99016 32070 99046 32122
rect 99046 32070 99058 32122
rect 99058 32070 99072 32122
rect 99096 32070 99110 32122
rect 99110 32070 99122 32122
rect 99122 32070 99152 32122
rect 99176 32070 99186 32122
rect 99186 32070 99232 32122
rect 98936 32068 98992 32070
rect 99016 32068 99072 32070
rect 99096 32068 99152 32070
rect 99176 32068 99232 32070
rect 98936 31034 98992 31036
rect 99016 31034 99072 31036
rect 99096 31034 99152 31036
rect 99176 31034 99232 31036
rect 98936 30982 98982 31034
rect 98982 30982 98992 31034
rect 99016 30982 99046 31034
rect 99046 30982 99058 31034
rect 99058 30982 99072 31034
rect 99096 30982 99110 31034
rect 99110 30982 99122 31034
rect 99122 30982 99152 31034
rect 99176 30982 99186 31034
rect 99186 30982 99232 31034
rect 98936 30980 98992 30982
rect 99016 30980 99072 30982
rect 99096 30980 99152 30982
rect 99176 30980 99232 30982
rect 99672 31578 99728 31580
rect 99752 31578 99808 31580
rect 99832 31578 99888 31580
rect 99912 31578 99968 31580
rect 99672 31526 99718 31578
rect 99718 31526 99728 31578
rect 99752 31526 99782 31578
rect 99782 31526 99794 31578
rect 99794 31526 99808 31578
rect 99832 31526 99846 31578
rect 99846 31526 99858 31578
rect 99858 31526 99888 31578
rect 99912 31526 99922 31578
rect 99922 31526 99968 31578
rect 99672 31524 99728 31526
rect 99752 31524 99808 31526
rect 99832 31524 99888 31526
rect 99912 31524 99968 31526
rect 98936 29946 98992 29948
rect 99016 29946 99072 29948
rect 99096 29946 99152 29948
rect 99176 29946 99232 29948
rect 98936 29894 98982 29946
rect 98982 29894 98992 29946
rect 99016 29894 99046 29946
rect 99046 29894 99058 29946
rect 99058 29894 99072 29946
rect 99096 29894 99110 29946
rect 99110 29894 99122 29946
rect 99122 29894 99152 29946
rect 99176 29894 99186 29946
rect 99186 29894 99232 29946
rect 98936 29892 98992 29894
rect 99016 29892 99072 29894
rect 99096 29892 99152 29894
rect 99176 29892 99232 29894
rect 98936 28858 98992 28860
rect 99016 28858 99072 28860
rect 99096 28858 99152 28860
rect 99176 28858 99232 28860
rect 98936 28806 98982 28858
rect 98982 28806 98992 28858
rect 99016 28806 99046 28858
rect 99046 28806 99058 28858
rect 99058 28806 99072 28858
rect 99096 28806 99110 28858
rect 99110 28806 99122 28858
rect 99122 28806 99152 28858
rect 99176 28806 99186 28858
rect 99186 28806 99232 28858
rect 98936 28804 98992 28806
rect 99016 28804 99072 28806
rect 99096 28804 99152 28806
rect 99176 28804 99232 28806
rect 98936 27770 98992 27772
rect 99016 27770 99072 27772
rect 99096 27770 99152 27772
rect 99176 27770 99232 27772
rect 98936 27718 98982 27770
rect 98982 27718 98992 27770
rect 99016 27718 99046 27770
rect 99046 27718 99058 27770
rect 99058 27718 99072 27770
rect 99096 27718 99110 27770
rect 99110 27718 99122 27770
rect 99122 27718 99152 27770
rect 99176 27718 99186 27770
rect 99186 27718 99232 27770
rect 98936 27716 98992 27718
rect 99016 27716 99072 27718
rect 99096 27716 99152 27718
rect 99176 27716 99232 27718
rect 98936 26682 98992 26684
rect 99016 26682 99072 26684
rect 99096 26682 99152 26684
rect 99176 26682 99232 26684
rect 98936 26630 98982 26682
rect 98982 26630 98992 26682
rect 99016 26630 99046 26682
rect 99046 26630 99058 26682
rect 99058 26630 99072 26682
rect 99096 26630 99110 26682
rect 99110 26630 99122 26682
rect 99122 26630 99152 26682
rect 99176 26630 99186 26682
rect 99186 26630 99232 26682
rect 98936 26628 98992 26630
rect 99016 26628 99072 26630
rect 99096 26628 99152 26630
rect 99176 26628 99232 26630
rect 99672 30490 99728 30492
rect 99752 30490 99808 30492
rect 99832 30490 99888 30492
rect 99912 30490 99968 30492
rect 99672 30438 99718 30490
rect 99718 30438 99728 30490
rect 99752 30438 99782 30490
rect 99782 30438 99794 30490
rect 99794 30438 99808 30490
rect 99832 30438 99846 30490
rect 99846 30438 99858 30490
rect 99858 30438 99888 30490
rect 99912 30438 99922 30490
rect 99922 30438 99968 30490
rect 99672 30436 99728 30438
rect 99752 30436 99808 30438
rect 99832 30436 99888 30438
rect 99912 30436 99968 30438
rect 99672 29402 99728 29404
rect 99752 29402 99808 29404
rect 99832 29402 99888 29404
rect 99912 29402 99968 29404
rect 99672 29350 99718 29402
rect 99718 29350 99728 29402
rect 99752 29350 99782 29402
rect 99782 29350 99794 29402
rect 99794 29350 99808 29402
rect 99832 29350 99846 29402
rect 99846 29350 99858 29402
rect 99858 29350 99888 29402
rect 99912 29350 99922 29402
rect 99922 29350 99968 29402
rect 99672 29348 99728 29350
rect 99752 29348 99808 29350
rect 99832 29348 99888 29350
rect 99912 29348 99968 29350
rect 99672 28314 99728 28316
rect 99752 28314 99808 28316
rect 99832 28314 99888 28316
rect 99912 28314 99968 28316
rect 99672 28262 99718 28314
rect 99718 28262 99728 28314
rect 99752 28262 99782 28314
rect 99782 28262 99794 28314
rect 99794 28262 99808 28314
rect 99832 28262 99846 28314
rect 99846 28262 99858 28314
rect 99858 28262 99888 28314
rect 99912 28262 99922 28314
rect 99922 28262 99968 28314
rect 99672 28260 99728 28262
rect 99752 28260 99808 28262
rect 99832 28260 99888 28262
rect 99912 28260 99968 28262
rect 99672 27226 99728 27228
rect 99752 27226 99808 27228
rect 99832 27226 99888 27228
rect 99912 27226 99968 27228
rect 99672 27174 99718 27226
rect 99718 27174 99728 27226
rect 99752 27174 99782 27226
rect 99782 27174 99794 27226
rect 99794 27174 99808 27226
rect 99832 27174 99846 27226
rect 99846 27174 99858 27226
rect 99858 27174 99888 27226
rect 99912 27174 99922 27226
rect 99922 27174 99968 27226
rect 99672 27172 99728 27174
rect 99752 27172 99808 27174
rect 99832 27172 99888 27174
rect 99912 27172 99968 27174
rect 99672 26138 99728 26140
rect 99752 26138 99808 26140
rect 99832 26138 99888 26140
rect 99912 26138 99968 26140
rect 99672 26086 99718 26138
rect 99718 26086 99728 26138
rect 99752 26086 99782 26138
rect 99782 26086 99794 26138
rect 99794 26086 99808 26138
rect 99832 26086 99846 26138
rect 99846 26086 99858 26138
rect 99858 26086 99888 26138
rect 99912 26086 99922 26138
rect 99922 26086 99968 26138
rect 99672 26084 99728 26086
rect 99752 26084 99808 26086
rect 99832 26084 99888 26086
rect 99912 26084 99968 26086
rect 98182 19080 98238 19136
rect 98936 25594 98992 25596
rect 99016 25594 99072 25596
rect 99096 25594 99152 25596
rect 99176 25594 99232 25596
rect 98936 25542 98982 25594
rect 98982 25542 98992 25594
rect 99016 25542 99046 25594
rect 99046 25542 99058 25594
rect 99058 25542 99072 25594
rect 99096 25542 99110 25594
rect 99110 25542 99122 25594
rect 99122 25542 99152 25594
rect 99176 25542 99186 25594
rect 99186 25542 99232 25594
rect 98936 25540 98992 25542
rect 99016 25540 99072 25542
rect 99096 25540 99152 25542
rect 99176 25540 99232 25542
rect 98936 24506 98992 24508
rect 99016 24506 99072 24508
rect 99096 24506 99152 24508
rect 99176 24506 99232 24508
rect 98936 24454 98982 24506
rect 98982 24454 98992 24506
rect 99016 24454 99046 24506
rect 99046 24454 99058 24506
rect 99058 24454 99072 24506
rect 99096 24454 99110 24506
rect 99110 24454 99122 24506
rect 99122 24454 99152 24506
rect 99176 24454 99186 24506
rect 99186 24454 99232 24506
rect 98936 24452 98992 24454
rect 99016 24452 99072 24454
rect 99096 24452 99152 24454
rect 99176 24452 99232 24454
rect 98936 23418 98992 23420
rect 99016 23418 99072 23420
rect 99096 23418 99152 23420
rect 99176 23418 99232 23420
rect 98936 23366 98982 23418
rect 98982 23366 98992 23418
rect 99016 23366 99046 23418
rect 99046 23366 99058 23418
rect 99058 23366 99072 23418
rect 99096 23366 99110 23418
rect 99110 23366 99122 23418
rect 99122 23366 99152 23418
rect 99176 23366 99186 23418
rect 99186 23366 99232 23418
rect 98936 23364 98992 23366
rect 99016 23364 99072 23366
rect 99096 23364 99152 23366
rect 99176 23364 99232 23366
rect 98936 22330 98992 22332
rect 99016 22330 99072 22332
rect 99096 22330 99152 22332
rect 99176 22330 99232 22332
rect 98936 22278 98982 22330
rect 98982 22278 98992 22330
rect 99016 22278 99046 22330
rect 99046 22278 99058 22330
rect 99058 22278 99072 22330
rect 99096 22278 99110 22330
rect 99110 22278 99122 22330
rect 99122 22278 99152 22330
rect 99176 22278 99186 22330
rect 99186 22278 99232 22330
rect 98936 22276 98992 22278
rect 99016 22276 99072 22278
rect 99096 22276 99152 22278
rect 99176 22276 99232 22278
rect 98936 21242 98992 21244
rect 99016 21242 99072 21244
rect 99096 21242 99152 21244
rect 99176 21242 99232 21244
rect 98936 21190 98982 21242
rect 98982 21190 98992 21242
rect 99016 21190 99046 21242
rect 99046 21190 99058 21242
rect 99058 21190 99072 21242
rect 99096 21190 99110 21242
rect 99110 21190 99122 21242
rect 99122 21190 99152 21242
rect 99176 21190 99186 21242
rect 99186 21190 99232 21242
rect 98936 21188 98992 21190
rect 99016 21188 99072 21190
rect 99096 21188 99152 21190
rect 99176 21188 99232 21190
rect 98936 20154 98992 20156
rect 99016 20154 99072 20156
rect 99096 20154 99152 20156
rect 99176 20154 99232 20156
rect 98936 20102 98982 20154
rect 98982 20102 98992 20154
rect 99016 20102 99046 20154
rect 99046 20102 99058 20154
rect 99058 20102 99072 20154
rect 99096 20102 99110 20154
rect 99110 20102 99122 20154
rect 99122 20102 99152 20154
rect 99176 20102 99186 20154
rect 99186 20102 99232 20154
rect 98936 20100 98992 20102
rect 99016 20100 99072 20102
rect 99096 20100 99152 20102
rect 99176 20100 99232 20102
rect 98936 19066 98992 19068
rect 99016 19066 99072 19068
rect 99096 19066 99152 19068
rect 99176 19066 99232 19068
rect 98936 19014 98982 19066
rect 98982 19014 98992 19066
rect 99016 19014 99046 19066
rect 99046 19014 99058 19066
rect 99058 19014 99072 19066
rect 99096 19014 99110 19066
rect 99110 19014 99122 19066
rect 99122 19014 99152 19066
rect 99176 19014 99186 19066
rect 99186 19014 99232 19066
rect 98936 19012 98992 19014
rect 99016 19012 99072 19014
rect 99096 19012 99152 19014
rect 99176 19012 99232 19014
rect 98936 17978 98992 17980
rect 99016 17978 99072 17980
rect 99096 17978 99152 17980
rect 99176 17978 99232 17980
rect 98936 17926 98982 17978
rect 98982 17926 98992 17978
rect 99016 17926 99046 17978
rect 99046 17926 99058 17978
rect 99058 17926 99072 17978
rect 99096 17926 99110 17978
rect 99110 17926 99122 17978
rect 99122 17926 99152 17978
rect 99176 17926 99186 17978
rect 99186 17926 99232 17978
rect 98936 17924 98992 17926
rect 99016 17924 99072 17926
rect 99096 17924 99152 17926
rect 99176 17924 99232 17926
rect 99672 25050 99728 25052
rect 99752 25050 99808 25052
rect 99832 25050 99888 25052
rect 99912 25050 99968 25052
rect 99672 24998 99718 25050
rect 99718 24998 99728 25050
rect 99752 24998 99782 25050
rect 99782 24998 99794 25050
rect 99794 24998 99808 25050
rect 99832 24998 99846 25050
rect 99846 24998 99858 25050
rect 99858 24998 99888 25050
rect 99912 24998 99922 25050
rect 99922 24998 99968 25050
rect 99672 24996 99728 24998
rect 99752 24996 99808 24998
rect 99832 24996 99888 24998
rect 99912 24996 99968 24998
rect 99672 23962 99728 23964
rect 99752 23962 99808 23964
rect 99832 23962 99888 23964
rect 99912 23962 99968 23964
rect 99672 23910 99718 23962
rect 99718 23910 99728 23962
rect 99752 23910 99782 23962
rect 99782 23910 99794 23962
rect 99794 23910 99808 23962
rect 99832 23910 99846 23962
rect 99846 23910 99858 23962
rect 99858 23910 99888 23962
rect 99912 23910 99922 23962
rect 99922 23910 99968 23962
rect 99672 23908 99728 23910
rect 99752 23908 99808 23910
rect 99832 23908 99888 23910
rect 99912 23908 99968 23910
rect 100482 25880 100538 25936
rect 99672 22874 99728 22876
rect 99752 22874 99808 22876
rect 99832 22874 99888 22876
rect 99912 22874 99968 22876
rect 99672 22822 99718 22874
rect 99718 22822 99728 22874
rect 99752 22822 99782 22874
rect 99782 22822 99794 22874
rect 99794 22822 99808 22874
rect 99832 22822 99846 22874
rect 99846 22822 99858 22874
rect 99858 22822 99888 22874
rect 99912 22822 99922 22874
rect 99922 22822 99968 22874
rect 99672 22820 99728 22822
rect 99752 22820 99808 22822
rect 99832 22820 99888 22822
rect 99912 22820 99968 22822
rect 99672 21786 99728 21788
rect 99752 21786 99808 21788
rect 99832 21786 99888 21788
rect 99912 21786 99968 21788
rect 99672 21734 99718 21786
rect 99718 21734 99728 21786
rect 99752 21734 99782 21786
rect 99782 21734 99794 21786
rect 99794 21734 99808 21786
rect 99832 21734 99846 21786
rect 99846 21734 99858 21786
rect 99858 21734 99888 21786
rect 99912 21734 99922 21786
rect 99922 21734 99968 21786
rect 99672 21732 99728 21734
rect 99752 21732 99808 21734
rect 99832 21732 99888 21734
rect 99912 21732 99968 21734
rect 99672 20698 99728 20700
rect 99752 20698 99808 20700
rect 99832 20698 99888 20700
rect 99912 20698 99968 20700
rect 99672 20646 99718 20698
rect 99718 20646 99728 20698
rect 99752 20646 99782 20698
rect 99782 20646 99794 20698
rect 99794 20646 99808 20698
rect 99832 20646 99846 20698
rect 99846 20646 99858 20698
rect 99858 20646 99888 20698
rect 99912 20646 99922 20698
rect 99922 20646 99968 20698
rect 99672 20644 99728 20646
rect 99752 20644 99808 20646
rect 99832 20644 99888 20646
rect 99912 20644 99968 20646
rect 99672 19610 99728 19612
rect 99752 19610 99808 19612
rect 99832 19610 99888 19612
rect 99912 19610 99968 19612
rect 99672 19558 99718 19610
rect 99718 19558 99728 19610
rect 99752 19558 99782 19610
rect 99782 19558 99794 19610
rect 99794 19558 99808 19610
rect 99832 19558 99846 19610
rect 99846 19558 99858 19610
rect 99858 19558 99888 19610
rect 99912 19558 99922 19610
rect 99922 19558 99968 19610
rect 99672 19556 99728 19558
rect 99752 19556 99808 19558
rect 99832 19556 99888 19558
rect 99912 19556 99968 19558
rect 99672 18522 99728 18524
rect 99752 18522 99808 18524
rect 99832 18522 99888 18524
rect 99912 18522 99968 18524
rect 99672 18470 99718 18522
rect 99718 18470 99728 18522
rect 99752 18470 99782 18522
rect 99782 18470 99794 18522
rect 99794 18470 99808 18522
rect 99832 18470 99846 18522
rect 99846 18470 99858 18522
rect 99858 18470 99888 18522
rect 99912 18470 99922 18522
rect 99922 18470 99968 18522
rect 99672 18468 99728 18470
rect 99752 18468 99808 18470
rect 99832 18468 99888 18470
rect 99912 18468 99968 18470
rect 99672 17434 99728 17436
rect 99752 17434 99808 17436
rect 99832 17434 99888 17436
rect 99912 17434 99968 17436
rect 99672 17382 99718 17434
rect 99718 17382 99728 17434
rect 99752 17382 99782 17434
rect 99782 17382 99794 17434
rect 99794 17382 99808 17434
rect 99832 17382 99846 17434
rect 99846 17382 99858 17434
rect 99858 17382 99888 17434
rect 99912 17382 99922 17434
rect 99922 17382 99968 17434
rect 99672 17380 99728 17382
rect 99752 17380 99808 17382
rect 99832 17380 99888 17382
rect 99912 17380 99968 17382
rect 99378 17312 99434 17368
rect 98936 16890 98992 16892
rect 99016 16890 99072 16892
rect 99096 16890 99152 16892
rect 99176 16890 99232 16892
rect 98936 16838 98982 16890
rect 98982 16838 98992 16890
rect 99016 16838 99046 16890
rect 99046 16838 99058 16890
rect 99058 16838 99072 16890
rect 99096 16838 99110 16890
rect 99110 16838 99122 16890
rect 99122 16838 99152 16890
rect 99176 16838 99186 16890
rect 99186 16838 99232 16890
rect 98936 16836 98992 16838
rect 99016 16836 99072 16838
rect 99096 16836 99152 16838
rect 99176 16836 99232 16838
rect 99672 16346 99728 16348
rect 99752 16346 99808 16348
rect 99832 16346 99888 16348
rect 99912 16346 99968 16348
rect 99672 16294 99718 16346
rect 99718 16294 99728 16346
rect 99752 16294 99782 16346
rect 99782 16294 99794 16346
rect 99794 16294 99808 16346
rect 99832 16294 99846 16346
rect 99846 16294 99858 16346
rect 99858 16294 99888 16346
rect 99912 16294 99922 16346
rect 99922 16294 99968 16346
rect 99672 16292 99728 16294
rect 99752 16292 99808 16294
rect 99832 16292 99888 16294
rect 99912 16292 99968 16294
rect 98550 16224 98606 16280
rect 98936 15802 98992 15804
rect 99016 15802 99072 15804
rect 99096 15802 99152 15804
rect 99176 15802 99232 15804
rect 98936 15750 98982 15802
rect 98982 15750 98992 15802
rect 99016 15750 99046 15802
rect 99046 15750 99058 15802
rect 99058 15750 99072 15802
rect 99096 15750 99110 15802
rect 99110 15750 99122 15802
rect 99122 15750 99152 15802
rect 99176 15750 99186 15802
rect 99186 15750 99232 15802
rect 98936 15748 98992 15750
rect 99016 15748 99072 15750
rect 99096 15748 99152 15750
rect 99176 15748 99232 15750
rect 99672 15258 99728 15260
rect 99752 15258 99808 15260
rect 99832 15258 99888 15260
rect 99912 15258 99968 15260
rect 99672 15206 99718 15258
rect 99718 15206 99728 15258
rect 99752 15206 99782 15258
rect 99782 15206 99794 15258
rect 99794 15206 99808 15258
rect 99832 15206 99846 15258
rect 99846 15206 99858 15258
rect 99858 15206 99888 15258
rect 99912 15206 99922 15258
rect 99922 15206 99968 15258
rect 99672 15204 99728 15206
rect 99752 15204 99808 15206
rect 99832 15204 99888 15206
rect 99912 15204 99968 15206
rect 98936 14714 98992 14716
rect 99016 14714 99072 14716
rect 99096 14714 99152 14716
rect 99176 14714 99232 14716
rect 98936 14662 98982 14714
rect 98982 14662 98992 14714
rect 99016 14662 99046 14714
rect 99046 14662 99058 14714
rect 99058 14662 99072 14714
rect 99096 14662 99110 14714
rect 99110 14662 99122 14714
rect 99122 14662 99152 14714
rect 99176 14662 99186 14714
rect 99186 14662 99232 14714
rect 98936 14660 98992 14662
rect 99016 14660 99072 14662
rect 99096 14660 99152 14662
rect 99176 14660 99232 14662
rect 99672 14170 99728 14172
rect 99752 14170 99808 14172
rect 99832 14170 99888 14172
rect 99912 14170 99968 14172
rect 99672 14118 99718 14170
rect 99718 14118 99728 14170
rect 99752 14118 99782 14170
rect 99782 14118 99794 14170
rect 99794 14118 99808 14170
rect 99832 14118 99846 14170
rect 99846 14118 99858 14170
rect 99858 14118 99888 14170
rect 99912 14118 99922 14170
rect 99922 14118 99968 14170
rect 99672 14116 99728 14118
rect 99752 14116 99808 14118
rect 99832 14116 99888 14118
rect 99912 14116 99968 14118
rect 98936 13626 98992 13628
rect 99016 13626 99072 13628
rect 99096 13626 99152 13628
rect 99176 13626 99232 13628
rect 98936 13574 98982 13626
rect 98982 13574 98992 13626
rect 99016 13574 99046 13626
rect 99046 13574 99058 13626
rect 99058 13574 99072 13626
rect 99096 13574 99110 13626
rect 99110 13574 99122 13626
rect 99122 13574 99152 13626
rect 99176 13574 99186 13626
rect 99186 13574 99232 13626
rect 98936 13572 98992 13574
rect 99016 13572 99072 13574
rect 99096 13572 99152 13574
rect 99176 13572 99232 13574
rect 99672 13082 99728 13084
rect 99752 13082 99808 13084
rect 99832 13082 99888 13084
rect 99912 13082 99968 13084
rect 99672 13030 99718 13082
rect 99718 13030 99728 13082
rect 99752 13030 99782 13082
rect 99782 13030 99794 13082
rect 99794 13030 99808 13082
rect 99832 13030 99846 13082
rect 99846 13030 99858 13082
rect 99858 13030 99888 13082
rect 99912 13030 99922 13082
rect 99922 13030 99968 13082
rect 99672 13028 99728 13030
rect 99752 13028 99808 13030
rect 99832 13028 99888 13030
rect 99912 13028 99968 13030
rect 98936 12538 98992 12540
rect 99016 12538 99072 12540
rect 99096 12538 99152 12540
rect 99176 12538 99232 12540
rect 98936 12486 98982 12538
rect 98982 12486 98992 12538
rect 99016 12486 99046 12538
rect 99046 12486 99058 12538
rect 99058 12486 99072 12538
rect 99096 12486 99110 12538
rect 99110 12486 99122 12538
rect 99122 12486 99152 12538
rect 99176 12486 99186 12538
rect 99186 12486 99232 12538
rect 98936 12484 98992 12486
rect 99016 12484 99072 12486
rect 99096 12484 99152 12486
rect 99176 12484 99232 12486
rect 99672 11994 99728 11996
rect 99752 11994 99808 11996
rect 99832 11994 99888 11996
rect 99912 11994 99968 11996
rect 99672 11942 99718 11994
rect 99718 11942 99728 11994
rect 99752 11942 99782 11994
rect 99782 11942 99794 11994
rect 99794 11942 99808 11994
rect 99832 11942 99846 11994
rect 99846 11942 99858 11994
rect 99858 11942 99888 11994
rect 99912 11942 99922 11994
rect 99922 11942 99968 11994
rect 99672 11940 99728 11942
rect 99752 11940 99808 11942
rect 99832 11940 99888 11942
rect 99912 11940 99968 11942
rect 98936 11450 98992 11452
rect 99016 11450 99072 11452
rect 99096 11450 99152 11452
rect 99176 11450 99232 11452
rect 98936 11398 98982 11450
rect 98982 11398 98992 11450
rect 99016 11398 99046 11450
rect 99046 11398 99058 11450
rect 99058 11398 99072 11450
rect 99096 11398 99110 11450
rect 99110 11398 99122 11450
rect 99122 11398 99152 11450
rect 99176 11398 99186 11450
rect 99186 11398 99232 11450
rect 98936 11396 98992 11398
rect 99016 11396 99072 11398
rect 99096 11396 99152 11398
rect 99176 11396 99232 11398
rect 99672 10906 99728 10908
rect 99752 10906 99808 10908
rect 99832 10906 99888 10908
rect 99912 10906 99968 10908
rect 99672 10854 99718 10906
rect 99718 10854 99728 10906
rect 99752 10854 99782 10906
rect 99782 10854 99794 10906
rect 99794 10854 99808 10906
rect 99832 10854 99846 10906
rect 99846 10854 99858 10906
rect 99858 10854 99888 10906
rect 99912 10854 99922 10906
rect 99922 10854 99968 10906
rect 99672 10852 99728 10854
rect 99752 10852 99808 10854
rect 99832 10852 99888 10854
rect 99912 10852 99968 10854
rect 98936 10362 98992 10364
rect 99016 10362 99072 10364
rect 99096 10362 99152 10364
rect 99176 10362 99232 10364
rect 98936 10310 98982 10362
rect 98982 10310 98992 10362
rect 99016 10310 99046 10362
rect 99046 10310 99058 10362
rect 99058 10310 99072 10362
rect 99096 10310 99110 10362
rect 99110 10310 99122 10362
rect 99122 10310 99152 10362
rect 99176 10310 99186 10362
rect 99186 10310 99232 10362
rect 98936 10308 98992 10310
rect 99016 10308 99072 10310
rect 99096 10308 99152 10310
rect 99176 10308 99232 10310
rect 99672 9818 99728 9820
rect 99752 9818 99808 9820
rect 99832 9818 99888 9820
rect 99912 9818 99968 9820
rect 99672 9766 99718 9818
rect 99718 9766 99728 9818
rect 99752 9766 99782 9818
rect 99782 9766 99794 9818
rect 99794 9766 99808 9818
rect 99832 9766 99846 9818
rect 99846 9766 99858 9818
rect 99858 9766 99888 9818
rect 99912 9766 99922 9818
rect 99922 9766 99968 9818
rect 99672 9764 99728 9766
rect 99752 9764 99808 9766
rect 99832 9764 99888 9766
rect 99912 9764 99968 9766
rect 98936 9274 98992 9276
rect 99016 9274 99072 9276
rect 99096 9274 99152 9276
rect 99176 9274 99232 9276
rect 98936 9222 98982 9274
rect 98982 9222 98992 9274
rect 99016 9222 99046 9274
rect 99046 9222 99058 9274
rect 99058 9222 99072 9274
rect 99096 9222 99110 9274
rect 99110 9222 99122 9274
rect 99122 9222 99152 9274
rect 99176 9222 99186 9274
rect 99186 9222 99232 9274
rect 98936 9220 98992 9222
rect 99016 9220 99072 9222
rect 99096 9220 99152 9222
rect 99176 9220 99232 9222
rect 99672 8730 99728 8732
rect 99752 8730 99808 8732
rect 99832 8730 99888 8732
rect 99912 8730 99968 8732
rect 99672 8678 99718 8730
rect 99718 8678 99728 8730
rect 99752 8678 99782 8730
rect 99782 8678 99794 8730
rect 99794 8678 99808 8730
rect 99832 8678 99846 8730
rect 99846 8678 99858 8730
rect 99858 8678 99888 8730
rect 99912 8678 99922 8730
rect 99922 8678 99968 8730
rect 99672 8676 99728 8678
rect 99752 8676 99808 8678
rect 99832 8676 99888 8678
rect 99912 8676 99968 8678
rect 98936 8186 98992 8188
rect 99016 8186 99072 8188
rect 99096 8186 99152 8188
rect 99176 8186 99232 8188
rect 98936 8134 98982 8186
rect 98982 8134 98992 8186
rect 99016 8134 99046 8186
rect 99046 8134 99058 8186
rect 99058 8134 99072 8186
rect 99096 8134 99110 8186
rect 99110 8134 99122 8186
rect 99122 8134 99152 8186
rect 99176 8134 99186 8186
rect 99186 8134 99232 8186
rect 98936 8132 98992 8134
rect 99016 8132 99072 8134
rect 99096 8132 99152 8134
rect 99176 8132 99232 8134
rect 99672 7642 99728 7644
rect 99752 7642 99808 7644
rect 99832 7642 99888 7644
rect 99912 7642 99968 7644
rect 99672 7590 99718 7642
rect 99718 7590 99728 7642
rect 99752 7590 99782 7642
rect 99782 7590 99794 7642
rect 99794 7590 99808 7642
rect 99832 7590 99846 7642
rect 99846 7590 99858 7642
rect 99858 7590 99888 7642
rect 99912 7590 99922 7642
rect 99922 7590 99968 7642
rect 99672 7588 99728 7590
rect 99752 7588 99808 7590
rect 99832 7588 99888 7590
rect 99912 7588 99968 7590
rect 98936 7098 98992 7100
rect 99016 7098 99072 7100
rect 99096 7098 99152 7100
rect 99176 7098 99232 7100
rect 98936 7046 98982 7098
rect 98982 7046 98992 7098
rect 99016 7046 99046 7098
rect 99046 7046 99058 7098
rect 99058 7046 99072 7098
rect 99096 7046 99110 7098
rect 99110 7046 99122 7098
rect 99122 7046 99152 7098
rect 99176 7046 99186 7098
rect 99186 7046 99232 7098
rect 98936 7044 98992 7046
rect 99016 7044 99072 7046
rect 99096 7044 99152 7046
rect 99176 7044 99232 7046
rect 99672 6554 99728 6556
rect 99752 6554 99808 6556
rect 99832 6554 99888 6556
rect 99912 6554 99968 6556
rect 99672 6502 99718 6554
rect 99718 6502 99728 6554
rect 99752 6502 99782 6554
rect 99782 6502 99794 6554
rect 99794 6502 99808 6554
rect 99832 6502 99846 6554
rect 99846 6502 99858 6554
rect 99858 6502 99888 6554
rect 99912 6502 99922 6554
rect 99922 6502 99968 6554
rect 99672 6500 99728 6502
rect 99752 6500 99808 6502
rect 99832 6500 99888 6502
rect 99912 6500 99968 6502
rect 98936 6010 98992 6012
rect 99016 6010 99072 6012
rect 99096 6010 99152 6012
rect 99176 6010 99232 6012
rect 98936 5958 98982 6010
rect 98982 5958 98992 6010
rect 99016 5958 99046 6010
rect 99046 5958 99058 6010
rect 99058 5958 99072 6010
rect 99096 5958 99110 6010
rect 99110 5958 99122 6010
rect 99122 5958 99152 6010
rect 99176 5958 99186 6010
rect 99186 5958 99232 6010
rect 98936 5956 98992 5958
rect 99016 5956 99072 5958
rect 99096 5956 99152 5958
rect 99176 5956 99232 5958
rect 99672 5466 99728 5468
rect 99752 5466 99808 5468
rect 99832 5466 99888 5468
rect 99912 5466 99968 5468
rect 99672 5414 99718 5466
rect 99718 5414 99728 5466
rect 99752 5414 99782 5466
rect 99782 5414 99794 5466
rect 99794 5414 99808 5466
rect 99832 5414 99846 5466
rect 99846 5414 99858 5466
rect 99858 5414 99888 5466
rect 99912 5414 99922 5466
rect 99922 5414 99968 5466
rect 99672 5412 99728 5414
rect 99752 5412 99808 5414
rect 99832 5412 99888 5414
rect 99912 5412 99968 5414
rect 98936 4922 98992 4924
rect 99016 4922 99072 4924
rect 99096 4922 99152 4924
rect 99176 4922 99232 4924
rect 98936 4870 98982 4922
rect 98982 4870 98992 4922
rect 99016 4870 99046 4922
rect 99046 4870 99058 4922
rect 99058 4870 99072 4922
rect 99096 4870 99110 4922
rect 99110 4870 99122 4922
rect 99122 4870 99152 4922
rect 99176 4870 99186 4922
rect 99186 4870 99232 4922
rect 98936 4868 98992 4870
rect 99016 4868 99072 4870
rect 99096 4868 99152 4870
rect 99176 4868 99232 4870
rect 99672 4378 99728 4380
rect 99752 4378 99808 4380
rect 99832 4378 99888 4380
rect 99912 4378 99968 4380
rect 99672 4326 99718 4378
rect 99718 4326 99728 4378
rect 99752 4326 99782 4378
rect 99782 4326 99794 4378
rect 99794 4326 99808 4378
rect 99832 4326 99846 4378
rect 99846 4326 99858 4378
rect 99858 4326 99888 4378
rect 99912 4326 99922 4378
rect 99922 4326 99968 4378
rect 99672 4324 99728 4326
rect 99752 4324 99808 4326
rect 99832 4324 99888 4326
rect 99912 4324 99968 4326
rect 97998 3848 98054 3904
rect 98936 3834 98992 3836
rect 99016 3834 99072 3836
rect 99096 3834 99152 3836
rect 99176 3834 99232 3836
rect 98936 3782 98982 3834
rect 98982 3782 98992 3834
rect 99016 3782 99046 3834
rect 99046 3782 99058 3834
rect 99058 3782 99072 3834
rect 99096 3782 99110 3834
rect 99110 3782 99122 3834
rect 99122 3782 99152 3834
rect 99176 3782 99186 3834
rect 99186 3782 99232 3834
rect 98936 3780 98992 3782
rect 99016 3780 99072 3782
rect 99096 3780 99152 3782
rect 99176 3780 99232 3782
rect 97538 3712 97594 3768
rect 97354 3576 97410 3632
rect 17406 3440 17462 3496
rect 19982 3440 20038 3496
rect 20626 3440 20682 3496
rect 21914 3440 21970 3496
rect 24490 3440 24546 3496
rect 25778 3440 25834 3496
rect 27066 3440 27122 3496
rect 27710 3440 27766 3496
rect 30286 3440 30342 3496
rect 33506 3440 33562 3496
rect 34794 3440 34850 3496
rect 1680 3290 1736 3292
rect 1760 3290 1816 3292
rect 1680 3238 1690 3290
rect 1690 3238 1736 3290
rect 1760 3238 1806 3290
rect 1806 3238 1816 3290
rect 1680 3236 1736 3238
rect 1760 3236 1816 3238
rect 1312 2746 1368 2748
rect 1392 2746 1448 2748
rect 1312 2694 1322 2746
rect 1322 2694 1368 2746
rect 1392 2694 1438 2746
rect 1438 2694 1448 2746
rect 1312 2692 1368 2694
rect 1392 2692 1448 2694
rect 1680 2202 1736 2204
rect 1760 2202 1816 2204
rect 1680 2150 1690 2202
rect 1690 2150 1736 2202
rect 1760 2150 1806 2202
rect 1806 2150 1816 2202
rect 1680 2148 1736 2150
rect 1760 2148 1816 2150
rect 18694 2760 18750 2816
rect 23202 2760 23258 2816
rect 28998 2760 29054 2816
rect 31574 2760 31630 2816
rect 32862 2760 32918 2816
rect 99672 3290 99728 3292
rect 99752 3290 99808 3292
rect 99832 3290 99888 3292
rect 99912 3290 99968 3292
rect 99672 3238 99718 3290
rect 99718 3238 99728 3290
rect 99752 3238 99782 3290
rect 99782 3238 99794 3290
rect 99794 3238 99808 3290
rect 99832 3238 99846 3290
rect 99846 3238 99858 3290
rect 99858 3238 99888 3290
rect 99912 3238 99922 3290
rect 99922 3238 99968 3290
rect 99672 3236 99728 3238
rect 99752 3236 99808 3238
rect 99832 3236 99888 3238
rect 99912 3236 99968 3238
rect 36082 2760 36138 2816
rect 37370 2760 37426 2816
rect 98936 2746 98992 2748
rect 99016 2746 99072 2748
rect 99096 2746 99152 2748
rect 99176 2746 99232 2748
rect 98936 2694 98982 2746
rect 98982 2694 98992 2746
rect 99016 2694 99046 2746
rect 99046 2694 99058 2746
rect 99058 2694 99072 2746
rect 99096 2694 99110 2746
rect 99110 2694 99122 2746
rect 99122 2694 99152 2746
rect 99176 2694 99186 2746
rect 99186 2694 99232 2746
rect 98936 2692 98992 2694
rect 99016 2692 99072 2694
rect 99096 2692 99152 2694
rect 99176 2692 99232 2694
rect 99672 2202 99728 2204
rect 99752 2202 99808 2204
rect 99832 2202 99888 2204
rect 99912 2202 99968 2204
rect 99672 2150 99718 2202
rect 99718 2150 99728 2202
rect 99752 2150 99782 2202
rect 99782 2150 99794 2202
rect 99794 2150 99808 2202
rect 99832 2150 99846 2202
rect 99846 2150 99858 2202
rect 99858 2150 99888 2202
rect 99912 2150 99922 2202
rect 99922 2150 99968 2202
rect 99672 2148 99728 2150
rect 99752 2148 99808 2150
rect 99832 2148 99888 2150
rect 99912 2148 99968 2150
<< metal3 >>
rect 4210 101760 4526 101761
rect 4210 101696 4216 101760
rect 4280 101696 4296 101760
rect 4360 101696 4376 101760
rect 4440 101696 4456 101760
rect 4520 101696 4526 101760
rect 4210 101695 4526 101696
rect 34930 101760 35246 101761
rect 34930 101696 34936 101760
rect 35000 101696 35016 101760
rect 35080 101696 35096 101760
rect 35160 101696 35176 101760
rect 35240 101696 35246 101760
rect 34930 101695 35246 101696
rect 65650 101760 65966 101761
rect 65650 101696 65656 101760
rect 65720 101696 65736 101760
rect 65800 101696 65816 101760
rect 65880 101696 65896 101760
rect 65960 101696 65966 101760
rect 65650 101695 65966 101696
rect 96370 101760 96686 101761
rect 96370 101696 96376 101760
rect 96440 101696 96456 101760
rect 96520 101696 96536 101760
rect 96600 101696 96616 101760
rect 96680 101696 96686 101760
rect 96370 101695 96686 101696
rect 4870 101216 5186 101217
rect 4870 101152 4876 101216
rect 4940 101152 4956 101216
rect 5020 101152 5036 101216
rect 5100 101152 5116 101216
rect 5180 101152 5186 101216
rect 4870 101151 5186 101152
rect 35590 101216 35906 101217
rect 35590 101152 35596 101216
rect 35660 101152 35676 101216
rect 35740 101152 35756 101216
rect 35820 101152 35836 101216
rect 35900 101152 35906 101216
rect 35590 101151 35906 101152
rect 66310 101216 66626 101217
rect 66310 101152 66316 101216
rect 66380 101152 66396 101216
rect 66460 101152 66476 101216
rect 66540 101152 66556 101216
rect 66620 101152 66626 101216
rect 66310 101151 66626 101152
rect 97030 101216 97346 101217
rect 97030 101152 97036 101216
rect 97100 101152 97116 101216
rect 97180 101152 97196 101216
rect 97260 101152 97276 101216
rect 97340 101152 97346 101216
rect 97030 101151 97346 101152
rect 4210 100672 4526 100673
rect 4210 100608 4216 100672
rect 4280 100608 4296 100672
rect 4360 100608 4376 100672
rect 4440 100608 4456 100672
rect 4520 100608 4526 100672
rect 4210 100607 4526 100608
rect 34930 100672 35246 100673
rect 34930 100608 34936 100672
rect 35000 100608 35016 100672
rect 35080 100608 35096 100672
rect 35160 100608 35176 100672
rect 35240 100608 35246 100672
rect 34930 100607 35246 100608
rect 65650 100672 65966 100673
rect 65650 100608 65656 100672
rect 65720 100608 65736 100672
rect 65800 100608 65816 100672
rect 65880 100608 65896 100672
rect 65960 100608 65966 100672
rect 65650 100607 65966 100608
rect 96370 100672 96686 100673
rect 96370 100608 96376 100672
rect 96440 100608 96456 100672
rect 96520 100608 96536 100672
rect 96600 100608 96616 100672
rect 96680 100608 96686 100672
rect 96370 100607 96686 100608
rect 4870 100128 5186 100129
rect 4870 100064 4876 100128
rect 4940 100064 4956 100128
rect 5020 100064 5036 100128
rect 5100 100064 5116 100128
rect 5180 100064 5186 100128
rect 4870 100063 5186 100064
rect 35590 100128 35906 100129
rect 35590 100064 35596 100128
rect 35660 100064 35676 100128
rect 35740 100064 35756 100128
rect 35820 100064 35836 100128
rect 35900 100064 35906 100128
rect 35590 100063 35906 100064
rect 66310 100128 66626 100129
rect 66310 100064 66316 100128
rect 66380 100064 66396 100128
rect 66460 100064 66476 100128
rect 66540 100064 66556 100128
rect 66620 100064 66626 100128
rect 66310 100063 66626 100064
rect 97030 100128 97346 100129
rect 97030 100064 97036 100128
rect 97100 100064 97116 100128
rect 97180 100064 97196 100128
rect 97260 100064 97276 100128
rect 97340 100064 97346 100128
rect 97030 100063 97346 100064
rect 4210 99584 4526 99585
rect 4210 99520 4216 99584
rect 4280 99520 4296 99584
rect 4360 99520 4376 99584
rect 4440 99520 4456 99584
rect 4520 99520 4526 99584
rect 4210 99519 4526 99520
rect 34930 99584 35246 99585
rect 34930 99520 34936 99584
rect 35000 99520 35016 99584
rect 35080 99520 35096 99584
rect 35160 99520 35176 99584
rect 35240 99520 35246 99584
rect 34930 99519 35246 99520
rect 65650 99584 65966 99585
rect 65650 99520 65656 99584
rect 65720 99520 65736 99584
rect 65800 99520 65816 99584
rect 65880 99520 65896 99584
rect 65960 99520 65966 99584
rect 65650 99519 65966 99520
rect 96370 99584 96686 99585
rect 96370 99520 96376 99584
rect 96440 99520 96456 99584
rect 96520 99520 96536 99584
rect 96600 99520 96616 99584
rect 96680 99520 96686 99584
rect 96370 99519 96686 99520
rect 4870 99040 5186 99041
rect 4870 98976 4876 99040
rect 4940 98976 4956 99040
rect 5020 98976 5036 99040
rect 5100 98976 5116 99040
rect 5180 98976 5186 99040
rect 4870 98975 5186 98976
rect 35590 99040 35906 99041
rect 35590 98976 35596 99040
rect 35660 98976 35676 99040
rect 35740 98976 35756 99040
rect 35820 98976 35836 99040
rect 35900 98976 35906 99040
rect 35590 98975 35906 98976
rect 66310 99040 66626 99041
rect 66310 98976 66316 99040
rect 66380 98976 66396 99040
rect 66460 98976 66476 99040
rect 66540 98976 66556 99040
rect 66620 98976 66626 99040
rect 66310 98975 66626 98976
rect 97030 99040 97346 99041
rect 97030 98976 97036 99040
rect 97100 98976 97116 99040
rect 97180 98976 97196 99040
rect 97260 98976 97276 99040
rect 97340 98976 97346 99040
rect 97030 98975 97346 98976
rect 4210 98496 4526 98497
rect 4210 98432 4216 98496
rect 4280 98432 4296 98496
rect 4360 98432 4376 98496
rect 4440 98432 4456 98496
rect 4520 98432 4526 98496
rect 4210 98431 4526 98432
rect 34930 98496 35246 98497
rect 34930 98432 34936 98496
rect 35000 98432 35016 98496
rect 35080 98432 35096 98496
rect 35160 98432 35176 98496
rect 35240 98432 35246 98496
rect 34930 98431 35246 98432
rect 65650 98496 65966 98497
rect 65650 98432 65656 98496
rect 65720 98432 65736 98496
rect 65800 98432 65816 98496
rect 65880 98432 65896 98496
rect 65960 98432 65966 98496
rect 65650 98431 65966 98432
rect 96370 98496 96686 98497
rect 96370 98432 96376 98496
rect 96440 98432 96456 98496
rect 96520 98432 96536 98496
rect 96600 98432 96616 98496
rect 96680 98432 96686 98496
rect 96370 98431 96686 98432
rect 4870 97952 5186 97953
rect 4870 97888 4876 97952
rect 4940 97888 4956 97952
rect 5020 97888 5036 97952
rect 5100 97888 5116 97952
rect 5180 97888 5186 97952
rect 4870 97887 5186 97888
rect 35590 97952 35906 97953
rect 35590 97888 35596 97952
rect 35660 97888 35676 97952
rect 35740 97888 35756 97952
rect 35820 97888 35836 97952
rect 35900 97888 35906 97952
rect 35590 97887 35906 97888
rect 66310 97952 66626 97953
rect 66310 97888 66316 97952
rect 66380 97888 66396 97952
rect 66460 97888 66476 97952
rect 66540 97888 66556 97952
rect 66620 97888 66626 97952
rect 66310 97887 66626 97888
rect 97030 97952 97346 97953
rect 97030 97888 97036 97952
rect 97100 97888 97116 97952
rect 97180 97888 97196 97952
rect 97260 97888 97276 97952
rect 97340 97888 97346 97952
rect 97030 97887 97346 97888
rect 4210 97408 4526 97409
rect 4210 97344 4216 97408
rect 4280 97344 4296 97408
rect 4360 97344 4376 97408
rect 4440 97344 4456 97408
rect 4520 97344 4526 97408
rect 4210 97343 4526 97344
rect 34930 97408 35246 97409
rect 34930 97344 34936 97408
rect 35000 97344 35016 97408
rect 35080 97344 35096 97408
rect 35160 97344 35176 97408
rect 35240 97344 35246 97408
rect 34930 97343 35246 97344
rect 65650 97408 65966 97409
rect 65650 97344 65656 97408
rect 65720 97344 65736 97408
rect 65800 97344 65816 97408
rect 65880 97344 65896 97408
rect 65960 97344 65966 97408
rect 65650 97343 65966 97344
rect 96370 97408 96686 97409
rect 96370 97344 96376 97408
rect 96440 97344 96456 97408
rect 96520 97344 96536 97408
rect 96600 97344 96616 97408
rect 96680 97344 96686 97408
rect 96370 97343 96686 97344
rect 4870 96864 5186 96865
rect 4870 96800 4876 96864
rect 4940 96800 4956 96864
rect 5020 96800 5036 96864
rect 5100 96800 5116 96864
rect 5180 96800 5186 96864
rect 4870 96799 5186 96800
rect 35590 96864 35906 96865
rect 35590 96800 35596 96864
rect 35660 96800 35676 96864
rect 35740 96800 35756 96864
rect 35820 96800 35836 96864
rect 35900 96800 35906 96864
rect 35590 96799 35906 96800
rect 66310 96864 66626 96865
rect 66310 96800 66316 96864
rect 66380 96800 66396 96864
rect 66460 96800 66476 96864
rect 66540 96800 66556 96864
rect 66620 96800 66626 96864
rect 66310 96799 66626 96800
rect 97030 96864 97346 96865
rect 97030 96800 97036 96864
rect 97100 96800 97116 96864
rect 97180 96800 97196 96864
rect 97260 96800 97276 96864
rect 97340 96800 97346 96864
rect 97030 96799 97346 96800
rect 4210 96320 4526 96321
rect 4210 96256 4216 96320
rect 4280 96256 4296 96320
rect 4360 96256 4376 96320
rect 4440 96256 4456 96320
rect 4520 96256 4526 96320
rect 4210 96255 4526 96256
rect 34930 96320 35246 96321
rect 34930 96256 34936 96320
rect 35000 96256 35016 96320
rect 35080 96256 35096 96320
rect 35160 96256 35176 96320
rect 35240 96256 35246 96320
rect 34930 96255 35246 96256
rect 65650 96320 65966 96321
rect 65650 96256 65656 96320
rect 65720 96256 65736 96320
rect 65800 96256 65816 96320
rect 65880 96256 65896 96320
rect 65960 96256 65966 96320
rect 65650 96255 65966 96256
rect 96370 96320 96686 96321
rect 96370 96256 96376 96320
rect 96440 96256 96456 96320
rect 96520 96256 96536 96320
rect 96600 96256 96616 96320
rect 96680 96256 96686 96320
rect 96370 96255 96686 96256
rect 4870 95776 5186 95777
rect 4870 95712 4876 95776
rect 4940 95712 4956 95776
rect 5020 95712 5036 95776
rect 5100 95712 5116 95776
rect 5180 95712 5186 95776
rect 4870 95711 5186 95712
rect 35590 95776 35906 95777
rect 35590 95712 35596 95776
rect 35660 95712 35676 95776
rect 35740 95712 35756 95776
rect 35820 95712 35836 95776
rect 35900 95712 35906 95776
rect 35590 95711 35906 95712
rect 66310 95776 66626 95777
rect 66310 95712 66316 95776
rect 66380 95712 66396 95776
rect 66460 95712 66476 95776
rect 66540 95712 66556 95776
rect 66620 95712 66626 95776
rect 66310 95711 66626 95712
rect 97030 95776 97346 95777
rect 97030 95712 97036 95776
rect 97100 95712 97116 95776
rect 97180 95712 97196 95776
rect 97260 95712 97276 95776
rect 97340 95712 97346 95776
rect 97030 95711 97346 95712
rect 4210 95232 4526 95233
rect 4210 95168 4216 95232
rect 4280 95168 4296 95232
rect 4360 95168 4376 95232
rect 4440 95168 4456 95232
rect 4520 95168 4526 95232
rect 4210 95167 4526 95168
rect 34930 95232 35246 95233
rect 34930 95168 34936 95232
rect 35000 95168 35016 95232
rect 35080 95168 35096 95232
rect 35160 95168 35176 95232
rect 35240 95168 35246 95232
rect 34930 95167 35246 95168
rect 65650 95232 65966 95233
rect 65650 95168 65656 95232
rect 65720 95168 65736 95232
rect 65800 95168 65816 95232
rect 65880 95168 65896 95232
rect 65960 95168 65966 95232
rect 65650 95167 65966 95168
rect 96370 95232 96686 95233
rect 96370 95168 96376 95232
rect 96440 95168 96456 95232
rect 96520 95168 96536 95232
rect 96600 95168 96616 95232
rect 96680 95168 96686 95232
rect 96370 95167 96686 95168
rect 4870 94688 5186 94689
rect 4870 94624 4876 94688
rect 4940 94624 4956 94688
rect 5020 94624 5036 94688
rect 5100 94624 5116 94688
rect 5180 94624 5186 94688
rect 4870 94623 5186 94624
rect 35590 94688 35906 94689
rect 35590 94624 35596 94688
rect 35660 94624 35676 94688
rect 35740 94624 35756 94688
rect 35820 94624 35836 94688
rect 35900 94624 35906 94688
rect 35590 94623 35906 94624
rect 66310 94688 66626 94689
rect 66310 94624 66316 94688
rect 66380 94624 66396 94688
rect 66460 94624 66476 94688
rect 66540 94624 66556 94688
rect 66620 94624 66626 94688
rect 66310 94623 66626 94624
rect 97030 94688 97346 94689
rect 97030 94624 97036 94688
rect 97100 94624 97116 94688
rect 97180 94624 97196 94688
rect 97260 94624 97276 94688
rect 97340 94624 97346 94688
rect 97030 94623 97346 94624
rect 4210 94144 4526 94145
rect 4210 94080 4216 94144
rect 4280 94080 4296 94144
rect 4360 94080 4376 94144
rect 4440 94080 4456 94144
rect 4520 94080 4526 94144
rect 4210 94079 4526 94080
rect 34930 94144 35246 94145
rect 34930 94080 34936 94144
rect 35000 94080 35016 94144
rect 35080 94080 35096 94144
rect 35160 94080 35176 94144
rect 35240 94080 35246 94144
rect 34930 94079 35246 94080
rect 65650 94144 65966 94145
rect 65650 94080 65656 94144
rect 65720 94080 65736 94144
rect 65800 94080 65816 94144
rect 65880 94080 65896 94144
rect 65960 94080 65966 94144
rect 65650 94079 65966 94080
rect 96370 94144 96686 94145
rect 96370 94080 96376 94144
rect 96440 94080 96456 94144
rect 96520 94080 96536 94144
rect 96600 94080 96616 94144
rect 96680 94080 96686 94144
rect 96370 94079 96686 94080
rect 4870 93600 5186 93601
rect 4870 93536 4876 93600
rect 4940 93536 4956 93600
rect 5020 93536 5036 93600
rect 5100 93536 5116 93600
rect 5180 93536 5186 93600
rect 4870 93535 5186 93536
rect 35590 93600 35906 93601
rect 35590 93536 35596 93600
rect 35660 93536 35676 93600
rect 35740 93536 35756 93600
rect 35820 93536 35836 93600
rect 35900 93536 35906 93600
rect 35590 93535 35906 93536
rect 66310 93600 66626 93601
rect 66310 93536 66316 93600
rect 66380 93536 66396 93600
rect 66460 93536 66476 93600
rect 66540 93536 66556 93600
rect 66620 93536 66626 93600
rect 66310 93535 66626 93536
rect 97030 93600 97346 93601
rect 97030 93536 97036 93600
rect 97100 93536 97116 93600
rect 97180 93536 97196 93600
rect 97260 93536 97276 93600
rect 97340 93536 97346 93600
rect 97030 93535 97346 93536
rect 4210 93056 4526 93057
rect 4210 92992 4216 93056
rect 4280 92992 4296 93056
rect 4360 92992 4376 93056
rect 4440 92992 4456 93056
rect 4520 92992 4526 93056
rect 4210 92991 4526 92992
rect 34930 93056 35246 93057
rect 34930 92992 34936 93056
rect 35000 92992 35016 93056
rect 35080 92992 35096 93056
rect 35160 92992 35176 93056
rect 35240 92992 35246 93056
rect 34930 92991 35246 92992
rect 65650 93056 65966 93057
rect 65650 92992 65656 93056
rect 65720 92992 65736 93056
rect 65800 92992 65816 93056
rect 65880 92992 65896 93056
rect 65960 92992 65966 93056
rect 65650 92991 65966 92992
rect 96370 93056 96686 93057
rect 96370 92992 96376 93056
rect 96440 92992 96456 93056
rect 96520 92992 96536 93056
rect 96600 92992 96616 93056
rect 96680 92992 96686 93056
rect 96370 92991 96686 92992
rect 4870 92512 5186 92513
rect 4870 92448 4876 92512
rect 4940 92448 4956 92512
rect 5020 92448 5036 92512
rect 5100 92448 5116 92512
rect 5180 92448 5186 92512
rect 4870 92447 5186 92448
rect 35590 92512 35906 92513
rect 35590 92448 35596 92512
rect 35660 92448 35676 92512
rect 35740 92448 35756 92512
rect 35820 92448 35836 92512
rect 35900 92448 35906 92512
rect 35590 92447 35906 92448
rect 66310 92512 66626 92513
rect 66310 92448 66316 92512
rect 66380 92448 66396 92512
rect 66460 92448 66476 92512
rect 66540 92448 66556 92512
rect 66620 92448 66626 92512
rect 66310 92447 66626 92448
rect 97030 92512 97346 92513
rect 97030 92448 97036 92512
rect 97100 92448 97116 92512
rect 97180 92448 97196 92512
rect 97260 92448 97276 92512
rect 97340 92448 97346 92512
rect 97030 92447 97346 92448
rect 4210 91968 4526 91969
rect 4210 91904 4216 91968
rect 4280 91904 4296 91968
rect 4360 91904 4376 91968
rect 4440 91904 4456 91968
rect 4520 91904 4526 91968
rect 4210 91903 4526 91904
rect 34930 91968 35246 91969
rect 34930 91904 34936 91968
rect 35000 91904 35016 91968
rect 35080 91904 35096 91968
rect 35160 91904 35176 91968
rect 35240 91904 35246 91968
rect 34930 91903 35246 91904
rect 65650 91968 65966 91969
rect 65650 91904 65656 91968
rect 65720 91904 65736 91968
rect 65800 91904 65816 91968
rect 65880 91904 65896 91968
rect 65960 91904 65966 91968
rect 65650 91903 65966 91904
rect 96370 91968 96686 91969
rect 96370 91904 96376 91968
rect 96440 91904 96456 91968
rect 96520 91904 96536 91968
rect 96600 91904 96616 91968
rect 96680 91904 96686 91968
rect 96370 91903 96686 91904
rect 4870 91424 5186 91425
rect 4870 91360 4876 91424
rect 4940 91360 4956 91424
rect 5020 91360 5036 91424
rect 5100 91360 5116 91424
rect 5180 91360 5186 91424
rect 4870 91359 5186 91360
rect 35590 91424 35906 91425
rect 35590 91360 35596 91424
rect 35660 91360 35676 91424
rect 35740 91360 35756 91424
rect 35820 91360 35836 91424
rect 35900 91360 35906 91424
rect 35590 91359 35906 91360
rect 66310 91424 66626 91425
rect 66310 91360 66316 91424
rect 66380 91360 66396 91424
rect 66460 91360 66476 91424
rect 66540 91360 66556 91424
rect 66620 91360 66626 91424
rect 66310 91359 66626 91360
rect 97030 91424 97346 91425
rect 97030 91360 97036 91424
rect 97100 91360 97116 91424
rect 97180 91360 97196 91424
rect 97260 91360 97276 91424
rect 97340 91360 97346 91424
rect 97030 91359 97346 91360
rect 4210 90880 4526 90881
rect 4210 90816 4216 90880
rect 4280 90816 4296 90880
rect 4360 90816 4376 90880
rect 4440 90816 4456 90880
rect 4520 90816 4526 90880
rect 4210 90815 4526 90816
rect 34930 90880 35246 90881
rect 34930 90816 34936 90880
rect 35000 90816 35016 90880
rect 35080 90816 35096 90880
rect 35160 90816 35176 90880
rect 35240 90816 35246 90880
rect 34930 90815 35246 90816
rect 65650 90880 65966 90881
rect 65650 90816 65656 90880
rect 65720 90816 65736 90880
rect 65800 90816 65816 90880
rect 65880 90816 65896 90880
rect 65960 90816 65966 90880
rect 65650 90815 65966 90816
rect 96370 90880 96686 90881
rect 96370 90816 96376 90880
rect 96440 90816 96456 90880
rect 96520 90816 96536 90880
rect 96600 90816 96616 90880
rect 96680 90816 96686 90880
rect 96370 90815 96686 90816
rect 4870 90336 5186 90337
rect 4870 90272 4876 90336
rect 4940 90272 4956 90336
rect 5020 90272 5036 90336
rect 5100 90272 5116 90336
rect 5180 90272 5186 90336
rect 4870 90271 5186 90272
rect 35590 90336 35906 90337
rect 35590 90272 35596 90336
rect 35660 90272 35676 90336
rect 35740 90272 35756 90336
rect 35820 90272 35836 90336
rect 35900 90272 35906 90336
rect 35590 90271 35906 90272
rect 66310 90336 66626 90337
rect 66310 90272 66316 90336
rect 66380 90272 66396 90336
rect 66460 90272 66476 90336
rect 66540 90272 66556 90336
rect 66620 90272 66626 90336
rect 66310 90271 66626 90272
rect 97030 90336 97346 90337
rect 97030 90272 97036 90336
rect 97100 90272 97116 90336
rect 97180 90272 97196 90336
rect 97260 90272 97276 90336
rect 97340 90272 97346 90336
rect 97030 90271 97346 90272
rect 4210 89792 4526 89793
rect 4210 89728 4216 89792
rect 4280 89728 4296 89792
rect 4360 89728 4376 89792
rect 4440 89728 4456 89792
rect 4520 89728 4526 89792
rect 4210 89727 4526 89728
rect 34930 89792 35246 89793
rect 34930 89728 34936 89792
rect 35000 89728 35016 89792
rect 35080 89728 35096 89792
rect 35160 89728 35176 89792
rect 35240 89728 35246 89792
rect 34930 89727 35246 89728
rect 65650 89792 65966 89793
rect 65650 89728 65656 89792
rect 65720 89728 65736 89792
rect 65800 89728 65816 89792
rect 65880 89728 65896 89792
rect 65960 89728 65966 89792
rect 65650 89727 65966 89728
rect 96370 89792 96686 89793
rect 96370 89728 96376 89792
rect 96440 89728 96456 89792
rect 96520 89728 96536 89792
rect 96600 89728 96616 89792
rect 96680 89728 96686 89792
rect 96370 89727 96686 89728
rect 4870 89248 5186 89249
rect 4870 89184 4876 89248
rect 4940 89184 4956 89248
rect 5020 89184 5036 89248
rect 5100 89184 5116 89248
rect 5180 89184 5186 89248
rect 4870 89183 5186 89184
rect 35590 89248 35906 89249
rect 35590 89184 35596 89248
rect 35660 89184 35676 89248
rect 35740 89184 35756 89248
rect 35820 89184 35836 89248
rect 35900 89184 35906 89248
rect 35590 89183 35906 89184
rect 66310 89248 66626 89249
rect 66310 89184 66316 89248
rect 66380 89184 66396 89248
rect 66460 89184 66476 89248
rect 66540 89184 66556 89248
rect 66620 89184 66626 89248
rect 66310 89183 66626 89184
rect 97030 89248 97346 89249
rect 97030 89184 97036 89248
rect 97100 89184 97116 89248
rect 97180 89184 97196 89248
rect 97260 89184 97276 89248
rect 97340 89184 97346 89248
rect 97030 89183 97346 89184
rect 4210 88704 4526 88705
rect 4210 88640 4216 88704
rect 4280 88640 4296 88704
rect 4360 88640 4376 88704
rect 4440 88640 4456 88704
rect 4520 88640 4526 88704
rect 4210 88639 4526 88640
rect 34930 88704 35246 88705
rect 34930 88640 34936 88704
rect 35000 88640 35016 88704
rect 35080 88640 35096 88704
rect 35160 88640 35176 88704
rect 35240 88640 35246 88704
rect 34930 88639 35246 88640
rect 65650 88704 65966 88705
rect 65650 88640 65656 88704
rect 65720 88640 65736 88704
rect 65800 88640 65816 88704
rect 65880 88640 65896 88704
rect 65960 88640 65966 88704
rect 65650 88639 65966 88640
rect 96370 88704 96686 88705
rect 96370 88640 96376 88704
rect 96440 88640 96456 88704
rect 96520 88640 96536 88704
rect 96600 88640 96616 88704
rect 96680 88640 96686 88704
rect 96370 88639 96686 88640
rect 4870 88160 5186 88161
rect 4870 88096 4876 88160
rect 4940 88096 4956 88160
rect 5020 88096 5036 88160
rect 5100 88096 5116 88160
rect 5180 88096 5186 88160
rect 4870 88095 5186 88096
rect 35590 88160 35906 88161
rect 35590 88096 35596 88160
rect 35660 88096 35676 88160
rect 35740 88096 35756 88160
rect 35820 88096 35836 88160
rect 35900 88096 35906 88160
rect 35590 88095 35906 88096
rect 66310 88160 66626 88161
rect 66310 88096 66316 88160
rect 66380 88096 66396 88160
rect 66460 88096 66476 88160
rect 66540 88096 66556 88160
rect 66620 88096 66626 88160
rect 66310 88095 66626 88096
rect 97030 88160 97346 88161
rect 97030 88096 97036 88160
rect 97100 88096 97116 88160
rect 97180 88096 97196 88160
rect 97260 88096 97276 88160
rect 97340 88096 97346 88160
rect 97030 88095 97346 88096
rect 4210 87616 4526 87617
rect 4210 87552 4216 87616
rect 4280 87552 4296 87616
rect 4360 87552 4376 87616
rect 4440 87552 4456 87616
rect 4520 87552 4526 87616
rect 4210 87551 4526 87552
rect 34930 87616 35246 87617
rect 34930 87552 34936 87616
rect 35000 87552 35016 87616
rect 35080 87552 35096 87616
rect 35160 87552 35176 87616
rect 35240 87552 35246 87616
rect 34930 87551 35246 87552
rect 65650 87616 65966 87617
rect 65650 87552 65656 87616
rect 65720 87552 65736 87616
rect 65800 87552 65816 87616
rect 65880 87552 65896 87616
rect 65960 87552 65966 87616
rect 65650 87551 65966 87552
rect 96370 87616 96686 87617
rect 96370 87552 96376 87616
rect 96440 87552 96456 87616
rect 96520 87552 96536 87616
rect 96600 87552 96616 87616
rect 96680 87552 96686 87616
rect 96370 87551 96686 87552
rect 4870 87072 5186 87073
rect 4870 87008 4876 87072
rect 4940 87008 4956 87072
rect 5020 87008 5036 87072
rect 5100 87008 5116 87072
rect 5180 87008 5186 87072
rect 4870 87007 5186 87008
rect 35590 87072 35906 87073
rect 35590 87008 35596 87072
rect 35660 87008 35676 87072
rect 35740 87008 35756 87072
rect 35820 87008 35836 87072
rect 35900 87008 35906 87072
rect 35590 87007 35906 87008
rect 66310 87072 66626 87073
rect 66310 87008 66316 87072
rect 66380 87008 66396 87072
rect 66460 87008 66476 87072
rect 66540 87008 66556 87072
rect 66620 87008 66626 87072
rect 66310 87007 66626 87008
rect 97030 87072 97346 87073
rect 97030 87008 97036 87072
rect 97100 87008 97116 87072
rect 97180 87008 97196 87072
rect 97260 87008 97276 87072
rect 97340 87008 97346 87072
rect 97030 87007 97346 87008
rect 4210 86528 4526 86529
rect 4210 86464 4216 86528
rect 4280 86464 4296 86528
rect 4360 86464 4376 86528
rect 4440 86464 4456 86528
rect 4520 86464 4526 86528
rect 4210 86463 4526 86464
rect 34930 86528 35246 86529
rect 34930 86464 34936 86528
rect 35000 86464 35016 86528
rect 35080 86464 35096 86528
rect 35160 86464 35176 86528
rect 35240 86464 35246 86528
rect 34930 86463 35246 86464
rect 65650 86528 65966 86529
rect 65650 86464 65656 86528
rect 65720 86464 65736 86528
rect 65800 86464 65816 86528
rect 65880 86464 65896 86528
rect 65960 86464 65966 86528
rect 65650 86463 65966 86464
rect 96370 86528 96686 86529
rect 96370 86464 96376 86528
rect 96440 86464 96456 86528
rect 96520 86464 96536 86528
rect 96600 86464 96616 86528
rect 96680 86464 96686 86528
rect 96370 86463 96686 86464
rect 4870 85984 5186 85985
rect 4870 85920 4876 85984
rect 4940 85920 4956 85984
rect 5020 85920 5036 85984
rect 5100 85920 5116 85984
rect 5180 85920 5186 85984
rect 4870 85919 5186 85920
rect 35590 85984 35906 85985
rect 35590 85920 35596 85984
rect 35660 85920 35676 85984
rect 35740 85920 35756 85984
rect 35820 85920 35836 85984
rect 35900 85920 35906 85984
rect 35590 85919 35906 85920
rect 66310 85984 66626 85985
rect 66310 85920 66316 85984
rect 66380 85920 66396 85984
rect 66460 85920 66476 85984
rect 66540 85920 66556 85984
rect 66620 85920 66626 85984
rect 66310 85919 66626 85920
rect 97030 85984 97346 85985
rect 97030 85920 97036 85984
rect 97100 85920 97116 85984
rect 97180 85920 97196 85984
rect 97260 85920 97276 85984
rect 97340 85920 97346 85984
rect 97030 85919 97346 85920
rect 4210 85440 4526 85441
rect 4210 85376 4216 85440
rect 4280 85376 4296 85440
rect 4360 85376 4376 85440
rect 4440 85376 4456 85440
rect 4520 85376 4526 85440
rect 4210 85375 4526 85376
rect 34930 85440 35246 85441
rect 34930 85376 34936 85440
rect 35000 85376 35016 85440
rect 35080 85376 35096 85440
rect 35160 85376 35176 85440
rect 35240 85376 35246 85440
rect 34930 85375 35246 85376
rect 65650 85440 65966 85441
rect 65650 85376 65656 85440
rect 65720 85376 65736 85440
rect 65800 85376 65816 85440
rect 65880 85376 65896 85440
rect 65960 85376 65966 85440
rect 65650 85375 65966 85376
rect 96370 85440 96686 85441
rect 96370 85376 96376 85440
rect 96440 85376 96456 85440
rect 96520 85376 96536 85440
rect 96600 85376 96616 85440
rect 96680 85376 96686 85440
rect 96370 85375 96686 85376
rect 4870 84896 5186 84897
rect 4870 84832 4876 84896
rect 4940 84832 4956 84896
rect 5020 84832 5036 84896
rect 5100 84832 5116 84896
rect 5180 84832 5186 84896
rect 4870 84831 5186 84832
rect 35590 84896 35906 84897
rect 35590 84832 35596 84896
rect 35660 84832 35676 84896
rect 35740 84832 35756 84896
rect 35820 84832 35836 84896
rect 35900 84832 35906 84896
rect 35590 84831 35906 84832
rect 66310 84896 66626 84897
rect 66310 84832 66316 84896
rect 66380 84832 66396 84896
rect 66460 84832 66476 84896
rect 66540 84832 66556 84896
rect 66620 84832 66626 84896
rect 66310 84831 66626 84832
rect 97030 84896 97346 84897
rect 97030 84832 97036 84896
rect 97100 84832 97116 84896
rect 97180 84832 97196 84896
rect 97260 84832 97276 84896
rect 97340 84832 97346 84896
rect 97030 84831 97346 84832
rect 4210 84352 4526 84353
rect 4210 84288 4216 84352
rect 4280 84288 4296 84352
rect 4360 84288 4376 84352
rect 4440 84288 4456 84352
rect 4520 84288 4526 84352
rect 4210 84287 4526 84288
rect 34930 84352 35246 84353
rect 34930 84288 34936 84352
rect 35000 84288 35016 84352
rect 35080 84288 35096 84352
rect 35160 84288 35176 84352
rect 35240 84288 35246 84352
rect 34930 84287 35246 84288
rect 65650 84352 65966 84353
rect 65650 84288 65656 84352
rect 65720 84288 65736 84352
rect 65800 84288 65816 84352
rect 65880 84288 65896 84352
rect 65960 84288 65966 84352
rect 65650 84287 65966 84288
rect 96370 84352 96686 84353
rect 96370 84288 96376 84352
rect 96440 84288 96456 84352
rect 96520 84288 96536 84352
rect 96600 84288 96616 84352
rect 96680 84288 96686 84352
rect 96370 84287 96686 84288
rect 4870 83808 5186 83809
rect 4870 83744 4876 83808
rect 4940 83744 4956 83808
rect 5020 83744 5036 83808
rect 5100 83744 5116 83808
rect 5180 83744 5186 83808
rect 4870 83743 5186 83744
rect 35590 83808 35906 83809
rect 35590 83744 35596 83808
rect 35660 83744 35676 83808
rect 35740 83744 35756 83808
rect 35820 83744 35836 83808
rect 35900 83744 35906 83808
rect 35590 83743 35906 83744
rect 66310 83808 66626 83809
rect 66310 83744 66316 83808
rect 66380 83744 66396 83808
rect 66460 83744 66476 83808
rect 66540 83744 66556 83808
rect 66620 83744 66626 83808
rect 66310 83743 66626 83744
rect 97030 83808 97346 83809
rect 97030 83744 97036 83808
rect 97100 83744 97116 83808
rect 97180 83744 97196 83808
rect 97260 83744 97276 83808
rect 97340 83744 97346 83808
rect 97030 83743 97346 83744
rect 4210 83264 4526 83265
rect 4210 83200 4216 83264
rect 4280 83200 4296 83264
rect 4360 83200 4376 83264
rect 4440 83200 4456 83264
rect 4520 83200 4526 83264
rect 4210 83199 4526 83200
rect 34930 83264 35246 83265
rect 34930 83200 34936 83264
rect 35000 83200 35016 83264
rect 35080 83200 35096 83264
rect 35160 83200 35176 83264
rect 35240 83200 35246 83264
rect 34930 83199 35246 83200
rect 65650 83264 65966 83265
rect 65650 83200 65656 83264
rect 65720 83200 65736 83264
rect 65800 83200 65816 83264
rect 65880 83200 65896 83264
rect 65960 83200 65966 83264
rect 65650 83199 65966 83200
rect 96370 83264 96686 83265
rect 96370 83200 96376 83264
rect 96440 83200 96456 83264
rect 96520 83200 96536 83264
rect 96600 83200 96616 83264
rect 96680 83200 96686 83264
rect 96370 83199 96686 83200
rect 4870 82720 5186 82721
rect 4870 82656 4876 82720
rect 4940 82656 4956 82720
rect 5020 82656 5036 82720
rect 5100 82656 5116 82720
rect 5180 82656 5186 82720
rect 4870 82655 5186 82656
rect 35590 82720 35906 82721
rect 35590 82656 35596 82720
rect 35660 82656 35676 82720
rect 35740 82656 35756 82720
rect 35820 82656 35836 82720
rect 35900 82656 35906 82720
rect 35590 82655 35906 82656
rect 66310 82720 66626 82721
rect 66310 82656 66316 82720
rect 66380 82656 66396 82720
rect 66460 82656 66476 82720
rect 66540 82656 66556 82720
rect 66620 82656 66626 82720
rect 66310 82655 66626 82656
rect 97030 82720 97346 82721
rect 97030 82656 97036 82720
rect 97100 82656 97116 82720
rect 97180 82656 97196 82720
rect 97260 82656 97276 82720
rect 97340 82656 97346 82720
rect 97030 82655 97346 82656
rect 4210 82176 4526 82177
rect 4210 82112 4216 82176
rect 4280 82112 4296 82176
rect 4360 82112 4376 82176
rect 4440 82112 4456 82176
rect 4520 82112 4526 82176
rect 4210 82111 4526 82112
rect 34930 82176 35246 82177
rect 34930 82112 34936 82176
rect 35000 82112 35016 82176
rect 35080 82112 35096 82176
rect 35160 82112 35176 82176
rect 35240 82112 35246 82176
rect 34930 82111 35246 82112
rect 65650 82176 65966 82177
rect 65650 82112 65656 82176
rect 65720 82112 65736 82176
rect 65800 82112 65816 82176
rect 65880 82112 65896 82176
rect 65960 82112 65966 82176
rect 65650 82111 65966 82112
rect 96370 82176 96686 82177
rect 96370 82112 96376 82176
rect 96440 82112 96456 82176
rect 96520 82112 96536 82176
rect 96600 82112 96616 82176
rect 96680 82112 96686 82176
rect 96370 82111 96686 82112
rect 4870 81632 5186 81633
rect 4870 81568 4876 81632
rect 4940 81568 4956 81632
rect 5020 81568 5036 81632
rect 5100 81568 5116 81632
rect 5180 81568 5186 81632
rect 4870 81567 5186 81568
rect 35590 81632 35906 81633
rect 35590 81568 35596 81632
rect 35660 81568 35676 81632
rect 35740 81568 35756 81632
rect 35820 81568 35836 81632
rect 35900 81568 35906 81632
rect 35590 81567 35906 81568
rect 66310 81632 66626 81633
rect 66310 81568 66316 81632
rect 66380 81568 66396 81632
rect 66460 81568 66476 81632
rect 66540 81568 66556 81632
rect 66620 81568 66626 81632
rect 66310 81567 66626 81568
rect 97030 81632 97346 81633
rect 97030 81568 97036 81632
rect 97100 81568 97116 81632
rect 97180 81568 97196 81632
rect 97260 81568 97276 81632
rect 97340 81568 97346 81632
rect 97030 81567 97346 81568
rect 4210 81088 4526 81089
rect 4210 81024 4216 81088
rect 4280 81024 4296 81088
rect 4360 81024 4376 81088
rect 4440 81024 4456 81088
rect 4520 81024 4526 81088
rect 4210 81023 4526 81024
rect 34930 81088 35246 81089
rect 34930 81024 34936 81088
rect 35000 81024 35016 81088
rect 35080 81024 35096 81088
rect 35160 81024 35176 81088
rect 35240 81024 35246 81088
rect 34930 81023 35246 81024
rect 65650 81088 65966 81089
rect 65650 81024 65656 81088
rect 65720 81024 65736 81088
rect 65800 81024 65816 81088
rect 65880 81024 65896 81088
rect 65960 81024 65966 81088
rect 65650 81023 65966 81024
rect 96370 81088 96686 81089
rect 96370 81024 96376 81088
rect 96440 81024 96456 81088
rect 96520 81024 96536 81088
rect 96600 81024 96616 81088
rect 96680 81024 96686 81088
rect 96370 81023 96686 81024
rect 4870 80544 5186 80545
rect 4870 80480 4876 80544
rect 4940 80480 4956 80544
rect 5020 80480 5036 80544
rect 5100 80480 5116 80544
rect 5180 80480 5186 80544
rect 4870 80479 5186 80480
rect 35590 80544 35906 80545
rect 35590 80480 35596 80544
rect 35660 80480 35676 80544
rect 35740 80480 35756 80544
rect 35820 80480 35836 80544
rect 35900 80480 35906 80544
rect 35590 80479 35906 80480
rect 66310 80544 66626 80545
rect 66310 80480 66316 80544
rect 66380 80480 66396 80544
rect 66460 80480 66476 80544
rect 66540 80480 66556 80544
rect 66620 80480 66626 80544
rect 66310 80479 66626 80480
rect 97030 80544 97346 80545
rect 97030 80480 97036 80544
rect 97100 80480 97116 80544
rect 97180 80480 97196 80544
rect 97260 80480 97276 80544
rect 97340 80480 97346 80544
rect 97030 80479 97346 80480
rect 4210 80000 4526 80001
rect 4210 79936 4216 80000
rect 4280 79936 4296 80000
rect 4360 79936 4376 80000
rect 4440 79936 4456 80000
rect 4520 79936 4526 80000
rect 4210 79935 4526 79936
rect 34930 80000 35246 80001
rect 34930 79936 34936 80000
rect 35000 79936 35016 80000
rect 35080 79936 35096 80000
rect 35160 79936 35176 80000
rect 35240 79936 35246 80000
rect 34930 79935 35246 79936
rect 65650 80000 65966 80001
rect 65650 79936 65656 80000
rect 65720 79936 65736 80000
rect 65800 79936 65816 80000
rect 65880 79936 65896 80000
rect 65960 79936 65966 80000
rect 65650 79935 65966 79936
rect 96370 80000 96686 80001
rect 96370 79936 96376 80000
rect 96440 79936 96456 80000
rect 96520 79936 96536 80000
rect 96600 79936 96616 80000
rect 96680 79936 96686 80000
rect 96370 79935 96686 79936
rect 4870 79456 5186 79457
rect 4870 79392 4876 79456
rect 4940 79392 4956 79456
rect 5020 79392 5036 79456
rect 5100 79392 5116 79456
rect 5180 79392 5186 79456
rect 4870 79391 5186 79392
rect 35590 79456 35906 79457
rect 35590 79392 35596 79456
rect 35660 79392 35676 79456
rect 35740 79392 35756 79456
rect 35820 79392 35836 79456
rect 35900 79392 35906 79456
rect 35590 79391 35906 79392
rect 66310 79456 66626 79457
rect 66310 79392 66316 79456
rect 66380 79392 66396 79456
rect 66460 79392 66476 79456
rect 66540 79392 66556 79456
rect 66620 79392 66626 79456
rect 66310 79391 66626 79392
rect 97030 79456 97346 79457
rect 97030 79392 97036 79456
rect 97100 79392 97116 79456
rect 97180 79392 97196 79456
rect 97260 79392 97276 79456
rect 97340 79392 97346 79456
rect 97030 79391 97346 79392
rect 4210 78912 4526 78913
rect 4210 78848 4216 78912
rect 4280 78848 4296 78912
rect 4360 78848 4376 78912
rect 4440 78848 4456 78912
rect 4520 78848 4526 78912
rect 4210 78847 4526 78848
rect 34930 78912 35246 78913
rect 34930 78848 34936 78912
rect 35000 78848 35016 78912
rect 35080 78848 35096 78912
rect 35160 78848 35176 78912
rect 35240 78848 35246 78912
rect 34930 78847 35246 78848
rect 65650 78912 65966 78913
rect 65650 78848 65656 78912
rect 65720 78848 65736 78912
rect 65800 78848 65816 78912
rect 65880 78848 65896 78912
rect 65960 78848 65966 78912
rect 65650 78847 65966 78848
rect 96370 78912 96686 78913
rect 96370 78848 96376 78912
rect 96440 78848 96456 78912
rect 96520 78848 96536 78912
rect 96600 78848 96616 78912
rect 96680 78848 96686 78912
rect 96370 78847 96686 78848
rect 4870 78368 5186 78369
rect 4870 78304 4876 78368
rect 4940 78304 4956 78368
rect 5020 78304 5036 78368
rect 5100 78304 5116 78368
rect 5180 78304 5186 78368
rect 4870 78303 5186 78304
rect 35590 78368 35906 78369
rect 35590 78304 35596 78368
rect 35660 78304 35676 78368
rect 35740 78304 35756 78368
rect 35820 78304 35836 78368
rect 35900 78304 35906 78368
rect 35590 78303 35906 78304
rect 66310 78368 66626 78369
rect 66310 78304 66316 78368
rect 66380 78304 66396 78368
rect 66460 78304 66476 78368
rect 66540 78304 66556 78368
rect 66620 78304 66626 78368
rect 66310 78303 66626 78304
rect 97030 78368 97346 78369
rect 97030 78304 97036 78368
rect 97100 78304 97116 78368
rect 97180 78304 97196 78368
rect 97260 78304 97276 78368
rect 97340 78304 97346 78368
rect 97030 78303 97346 78304
rect 4210 77824 4526 77825
rect 4210 77760 4216 77824
rect 4280 77760 4296 77824
rect 4360 77760 4376 77824
rect 4440 77760 4456 77824
rect 4520 77760 4526 77824
rect 4210 77759 4526 77760
rect 34930 77824 35246 77825
rect 34930 77760 34936 77824
rect 35000 77760 35016 77824
rect 35080 77760 35096 77824
rect 35160 77760 35176 77824
rect 35240 77760 35246 77824
rect 34930 77759 35246 77760
rect 65650 77824 65966 77825
rect 65650 77760 65656 77824
rect 65720 77760 65736 77824
rect 65800 77760 65816 77824
rect 65880 77760 65896 77824
rect 65960 77760 65966 77824
rect 65650 77759 65966 77760
rect 96370 77824 96686 77825
rect 96370 77760 96376 77824
rect 96440 77760 96456 77824
rect 96520 77760 96536 77824
rect 96600 77760 96616 77824
rect 96680 77760 96686 77824
rect 96370 77759 96686 77760
rect 4870 77280 5186 77281
rect 4870 77216 4876 77280
rect 4940 77216 4956 77280
rect 5020 77216 5036 77280
rect 5100 77216 5116 77280
rect 5180 77216 5186 77280
rect 4870 77215 5186 77216
rect 35590 77280 35906 77281
rect 35590 77216 35596 77280
rect 35660 77216 35676 77280
rect 35740 77216 35756 77280
rect 35820 77216 35836 77280
rect 35900 77216 35906 77280
rect 35590 77215 35906 77216
rect 66310 77280 66626 77281
rect 66310 77216 66316 77280
rect 66380 77216 66396 77280
rect 66460 77216 66476 77280
rect 66540 77216 66556 77280
rect 66620 77216 66626 77280
rect 66310 77215 66626 77216
rect 97030 77280 97346 77281
rect 97030 77216 97036 77280
rect 97100 77216 97116 77280
rect 97180 77216 97196 77280
rect 97260 77216 97276 77280
rect 97340 77216 97346 77280
rect 97030 77215 97346 77216
rect 45134 77012 45140 77076
rect 45204 77074 45210 77076
rect 49601 77074 49667 77077
rect 45204 77072 49667 77074
rect 45204 77016 49606 77072
rect 49662 77016 49667 77072
rect 45204 77014 49667 77016
rect 45204 77012 45210 77014
rect 49601 77011 49667 77014
rect 4210 76736 4526 76737
rect 4210 76672 4216 76736
rect 4280 76672 4296 76736
rect 4360 76672 4376 76736
rect 4440 76672 4456 76736
rect 4520 76672 4526 76736
rect 4210 76671 4526 76672
rect 34930 76736 35246 76737
rect 34930 76672 34936 76736
rect 35000 76672 35016 76736
rect 35080 76672 35096 76736
rect 35160 76672 35176 76736
rect 35240 76672 35246 76736
rect 34930 76671 35246 76672
rect 65650 76736 65966 76737
rect 65650 76672 65656 76736
rect 65720 76672 65736 76736
rect 65800 76672 65816 76736
rect 65880 76672 65896 76736
rect 65960 76672 65966 76736
rect 65650 76671 65966 76672
rect 96370 76736 96686 76737
rect 96370 76672 96376 76736
rect 96440 76672 96456 76736
rect 96520 76672 96536 76736
rect 96600 76672 96616 76736
rect 96680 76672 96686 76736
rect 96370 76671 96686 76672
rect 37590 76196 37596 76260
rect 37660 76258 37666 76260
rect 43621 76258 43687 76261
rect 37660 76256 43687 76258
rect 37660 76200 43626 76256
rect 43682 76200 43687 76256
rect 37660 76198 43687 76200
rect 37660 76196 37666 76198
rect 43621 76195 43687 76198
rect 4870 76192 5186 76193
rect 4870 76128 4876 76192
rect 4940 76128 4956 76192
rect 5020 76128 5036 76192
rect 5100 76128 5116 76192
rect 5180 76128 5186 76192
rect 4870 76127 5186 76128
rect 35590 76192 35906 76193
rect 35590 76128 35596 76192
rect 35660 76128 35676 76192
rect 35740 76128 35756 76192
rect 35820 76128 35836 76192
rect 35900 76128 35906 76192
rect 35590 76127 35906 76128
rect 66310 76192 66626 76193
rect 66310 76128 66316 76192
rect 66380 76128 66396 76192
rect 66460 76128 66476 76192
rect 66540 76128 66556 76192
rect 66620 76128 66626 76192
rect 66310 76127 66626 76128
rect 97030 76192 97346 76193
rect 97030 76128 97036 76192
rect 97100 76128 97116 76192
rect 97180 76128 97196 76192
rect 97260 76128 97276 76192
rect 97340 76128 97346 76192
rect 97030 76127 97346 76128
rect 42558 75924 42564 75988
rect 42628 75986 42634 75988
rect 47945 75986 48011 75989
rect 42628 75984 48011 75986
rect 42628 75928 47950 75984
rect 48006 75928 48011 75984
rect 42628 75926 48011 75928
rect 42628 75924 42634 75926
rect 47945 75923 48011 75926
rect 50102 75788 50108 75852
rect 50172 75850 50178 75852
rect 53281 75850 53347 75853
rect 50172 75848 53347 75850
rect 50172 75792 53286 75848
rect 53342 75792 53347 75848
rect 50172 75790 53347 75792
rect 50172 75788 50178 75790
rect 53281 75787 53347 75790
rect 4210 75648 4526 75649
rect 4210 75584 4216 75648
rect 4280 75584 4296 75648
rect 4360 75584 4376 75648
rect 4440 75584 4456 75648
rect 4520 75584 4526 75648
rect 4210 75583 4526 75584
rect 34930 75648 35246 75649
rect 34930 75584 34936 75648
rect 35000 75584 35016 75648
rect 35080 75584 35096 75648
rect 35160 75584 35176 75648
rect 35240 75584 35246 75648
rect 34930 75583 35246 75584
rect 65650 75648 65966 75649
rect 65650 75584 65656 75648
rect 65720 75584 65736 75648
rect 65800 75584 65816 75648
rect 65880 75584 65896 75648
rect 65960 75584 65966 75648
rect 65650 75583 65966 75584
rect 96370 75648 96686 75649
rect 96370 75584 96376 75648
rect 96440 75584 96456 75648
rect 96520 75584 96536 75648
rect 96600 75584 96616 75648
rect 96680 75584 96686 75648
rect 96370 75583 96686 75584
rect 4870 75104 5186 75105
rect 4870 75040 4876 75104
rect 4940 75040 4956 75104
rect 5020 75040 5036 75104
rect 5100 75040 5116 75104
rect 5180 75040 5186 75104
rect 4870 75039 5186 75040
rect 35590 75104 35906 75105
rect 35590 75040 35596 75104
rect 35660 75040 35676 75104
rect 35740 75040 35756 75104
rect 35820 75040 35836 75104
rect 35900 75040 35906 75104
rect 35590 75039 35906 75040
rect 66310 75104 66626 75105
rect 66310 75040 66316 75104
rect 66380 75040 66396 75104
rect 66460 75040 66476 75104
rect 66540 75040 66556 75104
rect 66620 75040 66626 75104
rect 66310 75039 66626 75040
rect 97030 75104 97346 75105
rect 97030 75040 97036 75104
rect 97100 75040 97116 75104
rect 97180 75040 97196 75104
rect 97260 75040 97276 75104
rect 97340 75040 97346 75104
rect 97030 75039 97346 75040
rect 40166 74564 40172 74628
rect 40236 74626 40242 74628
rect 45737 74626 45803 74629
rect 40236 74624 45803 74626
rect 40236 74568 45742 74624
rect 45798 74568 45803 74624
rect 40236 74566 45803 74568
rect 40236 74564 40242 74566
rect 45737 74563 45803 74566
rect 52494 74564 52500 74628
rect 52564 74626 52570 74628
rect 55581 74626 55647 74629
rect 52564 74624 55647 74626
rect 52564 74568 55586 74624
rect 55642 74568 55647 74624
rect 52564 74566 55647 74568
rect 52564 74564 52570 74566
rect 55581 74563 55647 74566
rect 4210 74560 4526 74561
rect 4210 74496 4216 74560
rect 4280 74496 4296 74560
rect 4360 74496 4376 74560
rect 4440 74496 4456 74560
rect 4520 74496 4526 74560
rect 4210 74495 4526 74496
rect 34930 74560 35246 74561
rect 34930 74496 34936 74560
rect 35000 74496 35016 74560
rect 35080 74496 35096 74560
rect 35160 74496 35176 74560
rect 35240 74496 35246 74560
rect 34930 74495 35246 74496
rect 65650 74560 65966 74561
rect 65650 74496 65656 74560
rect 65720 74496 65736 74560
rect 65800 74496 65816 74560
rect 65880 74496 65896 74560
rect 65960 74496 65966 74560
rect 65650 74495 65966 74496
rect 96370 74560 96686 74561
rect 96370 74496 96376 74560
rect 96440 74496 96456 74560
rect 96520 74496 96536 74560
rect 96600 74496 96616 74560
rect 96680 74496 96686 74560
rect 96370 74495 96686 74496
rect 4870 74016 5186 74017
rect 4870 73952 4876 74016
rect 4940 73952 4956 74016
rect 5020 73952 5036 74016
rect 5100 73952 5116 74016
rect 5180 73952 5186 74016
rect 4870 73951 5186 73952
rect 35590 74016 35906 74017
rect 35590 73952 35596 74016
rect 35660 73952 35676 74016
rect 35740 73952 35756 74016
rect 35820 73952 35836 74016
rect 35900 73952 35906 74016
rect 35590 73951 35906 73952
rect 66310 74016 66626 74017
rect 66310 73952 66316 74016
rect 66380 73952 66396 74016
rect 66460 73952 66476 74016
rect 66540 73952 66556 74016
rect 66620 73952 66626 74016
rect 66310 73951 66626 73952
rect 97030 74016 97346 74017
rect 97030 73952 97036 74016
rect 97100 73952 97116 74016
rect 97180 73952 97196 74016
rect 97260 73952 97276 74016
rect 97340 73952 97346 74016
rect 97030 73951 97346 73952
rect 55070 73884 55076 73948
rect 55140 73946 55146 73948
rect 57513 73946 57579 73949
rect 55140 73944 57579 73946
rect 55140 73888 57518 73944
rect 57574 73888 57579 73944
rect 55140 73886 57579 73888
rect 55140 73884 55146 73886
rect 57513 73883 57579 73886
rect 4210 73472 4526 73473
rect 4210 73408 4216 73472
rect 4280 73408 4296 73472
rect 4360 73408 4376 73472
rect 4440 73408 4456 73472
rect 4520 73408 4526 73472
rect 4210 73407 4526 73408
rect 34930 73472 35246 73473
rect 34930 73408 34936 73472
rect 35000 73408 35016 73472
rect 35080 73408 35096 73472
rect 35160 73408 35176 73472
rect 35240 73408 35246 73472
rect 34930 73407 35246 73408
rect 65650 73472 65966 73473
rect 65650 73408 65656 73472
rect 65720 73408 65736 73472
rect 65800 73408 65816 73472
rect 65880 73408 65896 73472
rect 65960 73408 65966 73472
rect 65650 73407 65966 73408
rect 96370 73472 96686 73473
rect 96370 73408 96376 73472
rect 96440 73408 96456 73472
rect 96520 73408 96536 73472
rect 96600 73408 96616 73472
rect 96680 73408 96686 73472
rect 96370 73407 96686 73408
rect 4870 72928 5186 72929
rect 4870 72864 4876 72928
rect 4940 72864 4956 72928
rect 5020 72864 5036 72928
rect 5100 72864 5116 72928
rect 5180 72864 5186 72928
rect 4870 72863 5186 72864
rect 35590 72928 35906 72929
rect 35590 72864 35596 72928
rect 35660 72864 35676 72928
rect 35740 72864 35756 72928
rect 35820 72864 35836 72928
rect 35900 72864 35906 72928
rect 35590 72863 35906 72864
rect 66310 72928 66626 72929
rect 66310 72864 66316 72928
rect 66380 72864 66396 72928
rect 66460 72864 66476 72928
rect 66540 72864 66556 72928
rect 66620 72864 66626 72928
rect 66310 72863 66626 72864
rect 97030 72928 97346 72929
rect 97030 72864 97036 72928
rect 97100 72864 97116 72928
rect 97180 72864 97196 72928
rect 97260 72864 97276 72928
rect 97340 72864 97346 72928
rect 97030 72863 97346 72864
rect 4210 72384 4526 72385
rect 4210 72320 4216 72384
rect 4280 72320 4296 72384
rect 4360 72320 4376 72384
rect 4440 72320 4456 72384
rect 4520 72320 4526 72384
rect 4210 72319 4526 72320
rect 34930 72384 35246 72385
rect 34930 72320 34936 72384
rect 35000 72320 35016 72384
rect 35080 72320 35096 72384
rect 35160 72320 35176 72384
rect 35240 72320 35246 72384
rect 34930 72319 35246 72320
rect 65650 72384 65966 72385
rect 65650 72320 65656 72384
rect 65720 72320 65736 72384
rect 65800 72320 65816 72384
rect 65880 72320 65896 72384
rect 65960 72320 65966 72384
rect 65650 72319 65966 72320
rect 96370 72384 96686 72385
rect 96370 72320 96376 72384
rect 96440 72320 96456 72384
rect 96520 72320 96536 72384
rect 96600 72320 96616 72384
rect 96680 72320 96686 72384
rect 96370 72319 96686 72320
rect 47526 71844 47532 71908
rect 47596 71906 47602 71908
rect 51257 71906 51323 71909
rect 47596 71904 51323 71906
rect 47596 71848 51262 71904
rect 51318 71848 51323 71904
rect 47596 71846 51323 71848
rect 47596 71844 47602 71846
rect 51257 71843 51323 71846
rect 4870 71840 5186 71841
rect 4870 71776 4876 71840
rect 4940 71776 4956 71840
rect 5020 71776 5036 71840
rect 5100 71776 5116 71840
rect 5180 71776 5186 71840
rect 4870 71775 5186 71776
rect 35590 71840 35906 71841
rect 35590 71776 35596 71840
rect 35660 71776 35676 71840
rect 35740 71776 35756 71840
rect 35820 71776 35836 71840
rect 35900 71776 35906 71840
rect 35590 71775 35906 71776
rect 66310 71840 66626 71841
rect 66310 71776 66316 71840
rect 66380 71776 66396 71840
rect 66460 71776 66476 71840
rect 66540 71776 66556 71840
rect 66620 71776 66626 71840
rect 66310 71775 66626 71776
rect 97030 71840 97346 71841
rect 97030 71776 97036 71840
rect 97100 71776 97116 71840
rect 97180 71776 97196 71840
rect 97260 71776 97276 71840
rect 97340 71776 97346 71840
rect 97030 71775 97346 71776
rect 4210 71296 4526 71297
rect 4210 71232 4216 71296
rect 4280 71232 4296 71296
rect 4360 71232 4376 71296
rect 4440 71232 4456 71296
rect 4520 71232 4526 71296
rect 4210 71231 4526 71232
rect 34930 71296 35246 71297
rect 34930 71232 34936 71296
rect 35000 71232 35016 71296
rect 35080 71232 35096 71296
rect 35160 71232 35176 71296
rect 35240 71232 35246 71296
rect 34930 71231 35246 71232
rect 65650 71296 65966 71297
rect 65650 71232 65656 71296
rect 65720 71232 65736 71296
rect 65800 71232 65816 71296
rect 65880 71232 65896 71296
rect 65960 71232 65966 71296
rect 65650 71231 65966 71232
rect 96370 71296 96686 71297
rect 96370 71232 96376 71296
rect 96440 71232 96456 71296
rect 96520 71232 96536 71296
rect 96600 71232 96616 71296
rect 96680 71232 96686 71296
rect 96370 71231 96686 71232
rect 4870 70752 5186 70753
rect 4870 70688 4876 70752
rect 4940 70688 4956 70752
rect 5020 70688 5036 70752
rect 5100 70688 5116 70752
rect 5180 70688 5186 70752
rect 4870 70687 5186 70688
rect 35590 70752 35906 70753
rect 35590 70688 35596 70752
rect 35660 70688 35676 70752
rect 35740 70688 35756 70752
rect 35820 70688 35836 70752
rect 35900 70688 35906 70752
rect 35590 70687 35906 70688
rect 66310 70752 66626 70753
rect 66310 70688 66316 70752
rect 66380 70688 66396 70752
rect 66460 70688 66476 70752
rect 66540 70688 66556 70752
rect 66620 70688 66626 70752
rect 66310 70687 66626 70688
rect 97030 70752 97346 70753
rect 97030 70688 97036 70752
rect 97100 70688 97116 70752
rect 97180 70688 97196 70752
rect 97260 70688 97276 70752
rect 97340 70688 97346 70752
rect 97030 70687 97346 70688
rect 4210 70208 4526 70209
rect 4210 70144 4216 70208
rect 4280 70144 4296 70208
rect 4360 70144 4376 70208
rect 4440 70144 4456 70208
rect 4520 70144 4526 70208
rect 4210 70143 4526 70144
rect 34930 70208 35246 70209
rect 34930 70144 34936 70208
rect 35000 70144 35016 70208
rect 35080 70144 35096 70208
rect 35160 70144 35176 70208
rect 35240 70144 35246 70208
rect 34930 70143 35246 70144
rect 65650 70208 65966 70209
rect 65650 70144 65656 70208
rect 65720 70144 65736 70208
rect 65800 70144 65816 70208
rect 65880 70144 65896 70208
rect 65960 70144 65966 70208
rect 65650 70143 65966 70144
rect 96370 70208 96686 70209
rect 96370 70144 96376 70208
rect 96440 70144 96456 70208
rect 96520 70144 96536 70208
rect 96600 70144 96616 70208
rect 96680 70144 96686 70208
rect 96370 70143 96686 70144
rect 4870 69664 5186 69665
rect 4870 69600 4876 69664
rect 4940 69600 4956 69664
rect 5020 69600 5036 69664
rect 5100 69600 5116 69664
rect 5180 69600 5186 69664
rect 4870 69599 5186 69600
rect 35590 69664 35906 69665
rect 35590 69600 35596 69664
rect 35660 69600 35676 69664
rect 35740 69600 35756 69664
rect 35820 69600 35836 69664
rect 35900 69600 35906 69664
rect 35590 69599 35906 69600
rect 66310 69664 66626 69665
rect 66310 69600 66316 69664
rect 66380 69600 66396 69664
rect 66460 69600 66476 69664
rect 66540 69600 66556 69664
rect 66620 69600 66626 69664
rect 66310 69599 66626 69600
rect 97030 69664 97346 69665
rect 97030 69600 97036 69664
rect 97100 69600 97116 69664
rect 97180 69600 97196 69664
rect 97260 69600 97276 69664
rect 97340 69600 97346 69664
rect 97030 69599 97346 69600
rect 4210 69120 4526 69121
rect 4210 69056 4216 69120
rect 4280 69056 4296 69120
rect 4360 69056 4376 69120
rect 4440 69056 4456 69120
rect 4520 69056 4526 69120
rect 4210 69055 4526 69056
rect 34930 69120 35246 69121
rect 34930 69056 34936 69120
rect 35000 69056 35016 69120
rect 35080 69056 35096 69120
rect 35160 69056 35176 69120
rect 35240 69056 35246 69120
rect 34930 69055 35246 69056
rect 65650 69120 65966 69121
rect 65650 69056 65656 69120
rect 65720 69056 65736 69120
rect 65800 69056 65816 69120
rect 65880 69056 65896 69120
rect 65960 69056 65966 69120
rect 65650 69055 65966 69056
rect 96370 69120 96686 69121
rect 96370 69056 96376 69120
rect 96440 69056 96456 69120
rect 96520 69056 96536 69120
rect 96600 69056 96616 69120
rect 96680 69056 96686 69120
rect 96370 69055 96686 69056
rect 4870 68576 5186 68577
rect 4870 68512 4876 68576
rect 4940 68512 4956 68576
rect 5020 68512 5036 68576
rect 5100 68512 5116 68576
rect 5180 68512 5186 68576
rect 4870 68511 5186 68512
rect 35590 68576 35906 68577
rect 35590 68512 35596 68576
rect 35660 68512 35676 68576
rect 35740 68512 35756 68576
rect 35820 68512 35836 68576
rect 35900 68512 35906 68576
rect 35590 68511 35906 68512
rect 66310 68576 66626 68577
rect 66310 68512 66316 68576
rect 66380 68512 66396 68576
rect 66460 68512 66476 68576
rect 66540 68512 66556 68576
rect 66620 68512 66626 68576
rect 66310 68511 66626 68512
rect 97030 68576 97346 68577
rect 97030 68512 97036 68576
rect 97100 68512 97116 68576
rect 97180 68512 97196 68576
rect 97260 68512 97276 68576
rect 97340 68512 97346 68576
rect 97030 68511 97346 68512
rect 4210 68032 4526 68033
rect 4210 67968 4216 68032
rect 4280 67968 4296 68032
rect 4360 67968 4376 68032
rect 4440 67968 4456 68032
rect 4520 67968 4526 68032
rect 4210 67967 4526 67968
rect 34930 68032 35246 68033
rect 34930 67968 34936 68032
rect 35000 67968 35016 68032
rect 35080 67968 35096 68032
rect 35160 67968 35176 68032
rect 35240 67968 35246 68032
rect 34930 67967 35246 67968
rect 65650 68032 65966 68033
rect 65650 67968 65656 68032
rect 65720 67968 65736 68032
rect 65800 67968 65816 68032
rect 65880 67968 65896 68032
rect 65960 67968 65966 68032
rect 65650 67967 65966 67968
rect 96370 68032 96686 68033
rect 96370 67968 96376 68032
rect 96440 67968 96456 68032
rect 96520 67968 96536 68032
rect 96600 67968 96616 68032
rect 96680 67968 96686 68032
rect 96370 67967 96686 67968
rect 4870 67488 5186 67489
rect 4870 67424 4876 67488
rect 4940 67424 4956 67488
rect 5020 67424 5036 67488
rect 5100 67424 5116 67488
rect 5180 67424 5186 67488
rect 4870 67423 5186 67424
rect 35590 67488 35906 67489
rect 35590 67424 35596 67488
rect 35660 67424 35676 67488
rect 35740 67424 35756 67488
rect 35820 67424 35836 67488
rect 35900 67424 35906 67488
rect 35590 67423 35906 67424
rect 66310 67488 66626 67489
rect 66310 67424 66316 67488
rect 66380 67424 66396 67488
rect 66460 67424 66476 67488
rect 66540 67424 66556 67488
rect 66620 67424 66626 67488
rect 66310 67423 66626 67424
rect 97030 67488 97346 67489
rect 97030 67424 97036 67488
rect 97100 67424 97116 67488
rect 97180 67424 97196 67488
rect 97260 67424 97276 67488
rect 97340 67424 97346 67488
rect 97030 67423 97346 67424
rect 4210 66944 4526 66945
rect 4210 66880 4216 66944
rect 4280 66880 4296 66944
rect 4360 66880 4376 66944
rect 4440 66880 4456 66944
rect 4520 66880 4526 66944
rect 4210 66879 4526 66880
rect 34930 66944 35246 66945
rect 34930 66880 34936 66944
rect 35000 66880 35016 66944
rect 35080 66880 35096 66944
rect 35160 66880 35176 66944
rect 35240 66880 35246 66944
rect 34930 66879 35246 66880
rect 65650 66944 65966 66945
rect 65650 66880 65656 66944
rect 65720 66880 65736 66944
rect 65800 66880 65816 66944
rect 65880 66880 65896 66944
rect 65960 66880 65966 66944
rect 65650 66879 65966 66880
rect 96370 66944 96686 66945
rect 96370 66880 96376 66944
rect 96440 66880 96456 66944
rect 96520 66880 96536 66944
rect 96600 66880 96616 66944
rect 96680 66880 96686 66944
rect 96370 66879 96686 66880
rect 4870 66400 5186 66401
rect 4870 66336 4876 66400
rect 4940 66336 4956 66400
rect 5020 66336 5036 66400
rect 5100 66336 5116 66400
rect 5180 66336 5186 66400
rect 4870 66335 5186 66336
rect 35590 66400 35906 66401
rect 35590 66336 35596 66400
rect 35660 66336 35676 66400
rect 35740 66336 35756 66400
rect 35820 66336 35836 66400
rect 35900 66336 35906 66400
rect 35590 66335 35906 66336
rect 66310 66400 66626 66401
rect 66310 66336 66316 66400
rect 66380 66336 66396 66400
rect 66460 66336 66476 66400
rect 66540 66336 66556 66400
rect 66620 66336 66626 66400
rect 66310 66335 66626 66336
rect 97030 66400 97346 66401
rect 97030 66336 97036 66400
rect 97100 66336 97116 66400
rect 97180 66336 97196 66400
rect 97260 66336 97276 66400
rect 97340 66336 97346 66400
rect 97030 66335 97346 66336
rect 4210 65856 4526 65857
rect 4210 65792 4216 65856
rect 4280 65792 4296 65856
rect 4360 65792 4376 65856
rect 4440 65792 4456 65856
rect 4520 65792 4526 65856
rect 4210 65791 4526 65792
rect 34930 65856 35246 65857
rect 34930 65792 34936 65856
rect 35000 65792 35016 65856
rect 35080 65792 35096 65856
rect 35160 65792 35176 65856
rect 35240 65792 35246 65856
rect 34930 65791 35246 65792
rect 65650 65856 65966 65857
rect 65650 65792 65656 65856
rect 65720 65792 65736 65856
rect 65800 65792 65816 65856
rect 65880 65792 65896 65856
rect 65960 65792 65966 65856
rect 65650 65791 65966 65792
rect 96370 65856 96686 65857
rect 96370 65792 96376 65856
rect 96440 65792 96456 65856
rect 96520 65792 96536 65856
rect 96600 65792 96616 65856
rect 96680 65792 96686 65856
rect 96370 65791 96686 65792
rect 4870 65312 5186 65313
rect 4870 65248 4876 65312
rect 4940 65248 4956 65312
rect 5020 65248 5036 65312
rect 5100 65248 5116 65312
rect 5180 65248 5186 65312
rect 4870 65247 5186 65248
rect 35590 65312 35906 65313
rect 35590 65248 35596 65312
rect 35660 65248 35676 65312
rect 35740 65248 35756 65312
rect 35820 65248 35836 65312
rect 35900 65248 35906 65312
rect 35590 65247 35906 65248
rect 66310 65312 66626 65313
rect 66310 65248 66316 65312
rect 66380 65248 66396 65312
rect 66460 65248 66476 65312
rect 66540 65248 66556 65312
rect 66620 65248 66626 65312
rect 66310 65247 66626 65248
rect 97030 65312 97346 65313
rect 97030 65248 97036 65312
rect 97100 65248 97116 65312
rect 97180 65248 97196 65312
rect 97260 65248 97276 65312
rect 97340 65248 97346 65312
rect 97030 65247 97346 65248
rect 4210 64768 4526 64769
rect 4210 64704 4216 64768
rect 4280 64704 4296 64768
rect 4360 64704 4376 64768
rect 4440 64704 4456 64768
rect 4520 64704 4526 64768
rect 4210 64703 4526 64704
rect 34930 64768 35246 64769
rect 34930 64704 34936 64768
rect 35000 64704 35016 64768
rect 35080 64704 35096 64768
rect 35160 64704 35176 64768
rect 35240 64704 35246 64768
rect 34930 64703 35246 64704
rect 65650 64768 65966 64769
rect 65650 64704 65656 64768
rect 65720 64704 65736 64768
rect 65800 64704 65816 64768
rect 65880 64704 65896 64768
rect 65960 64704 65966 64768
rect 65650 64703 65966 64704
rect 96370 64768 96686 64769
rect 96370 64704 96376 64768
rect 96440 64704 96456 64768
rect 96520 64704 96536 64768
rect 96600 64704 96616 64768
rect 96680 64704 96686 64768
rect 96370 64703 96686 64704
rect 4870 64224 5186 64225
rect 4870 64160 4876 64224
rect 4940 64160 4956 64224
rect 5020 64160 5036 64224
rect 5100 64160 5116 64224
rect 5180 64160 5186 64224
rect 4870 64159 5186 64160
rect 35590 64224 35906 64225
rect 35590 64160 35596 64224
rect 35660 64160 35676 64224
rect 35740 64160 35756 64224
rect 35820 64160 35836 64224
rect 35900 64160 35906 64224
rect 35590 64159 35906 64160
rect 66310 64224 66626 64225
rect 66310 64160 66316 64224
rect 66380 64160 66396 64224
rect 66460 64160 66476 64224
rect 66540 64160 66556 64224
rect 66620 64160 66626 64224
rect 66310 64159 66626 64160
rect 97030 64224 97346 64225
rect 97030 64160 97036 64224
rect 97100 64160 97116 64224
rect 97180 64160 97196 64224
rect 97260 64160 97276 64224
rect 97340 64160 97346 64224
rect 97030 64159 97346 64160
rect 4210 63680 4526 63681
rect 4210 63616 4216 63680
rect 4280 63616 4296 63680
rect 4360 63616 4376 63680
rect 4440 63616 4456 63680
rect 4520 63616 4526 63680
rect 4210 63615 4526 63616
rect 34930 63680 35246 63681
rect 34930 63616 34936 63680
rect 35000 63616 35016 63680
rect 35080 63616 35096 63680
rect 35160 63616 35176 63680
rect 35240 63616 35246 63680
rect 34930 63615 35246 63616
rect 65650 63680 65966 63681
rect 65650 63616 65656 63680
rect 65720 63616 65736 63680
rect 65800 63616 65816 63680
rect 65880 63616 65896 63680
rect 65960 63616 65966 63680
rect 65650 63615 65966 63616
rect 96370 63680 96686 63681
rect 96370 63616 96376 63680
rect 96440 63616 96456 63680
rect 96520 63616 96536 63680
rect 96600 63616 96616 63680
rect 96680 63616 96686 63680
rect 96370 63615 96686 63616
rect 4870 63136 5186 63137
rect 4870 63072 4876 63136
rect 4940 63072 4956 63136
rect 5020 63072 5036 63136
rect 5100 63072 5116 63136
rect 5180 63072 5186 63136
rect 4870 63071 5186 63072
rect 35590 63136 35906 63137
rect 35590 63072 35596 63136
rect 35660 63072 35676 63136
rect 35740 63072 35756 63136
rect 35820 63072 35836 63136
rect 35900 63072 35906 63136
rect 35590 63071 35906 63072
rect 66310 63136 66626 63137
rect 66310 63072 66316 63136
rect 66380 63072 66396 63136
rect 66460 63072 66476 63136
rect 66540 63072 66556 63136
rect 66620 63072 66626 63136
rect 66310 63071 66626 63072
rect 97030 63136 97346 63137
rect 97030 63072 97036 63136
rect 97100 63072 97116 63136
rect 97180 63072 97196 63136
rect 97260 63072 97276 63136
rect 97340 63072 97346 63136
rect 97030 63071 97346 63072
rect 35382 62732 35388 62796
rect 35452 62794 35458 62796
rect 41781 62794 41847 62797
rect 35452 62792 41847 62794
rect 35452 62736 41786 62792
rect 41842 62736 41847 62792
rect 35452 62734 41847 62736
rect 35452 62732 35458 62734
rect 41781 62731 41847 62734
rect 100385 62658 100451 62661
rect 101162 62658 101962 62688
rect 100385 62656 101962 62658
rect 100385 62600 100390 62656
rect 100446 62600 101962 62656
rect 100385 62598 101962 62600
rect 100385 62595 100451 62598
rect 4210 62592 4526 62593
rect 4210 62528 4216 62592
rect 4280 62528 4296 62592
rect 4360 62528 4376 62592
rect 4440 62528 4456 62592
rect 4520 62528 4526 62592
rect 4210 62527 4526 62528
rect 34930 62592 35246 62593
rect 34930 62528 34936 62592
rect 35000 62528 35016 62592
rect 35080 62528 35096 62592
rect 35160 62528 35176 62592
rect 35240 62528 35246 62592
rect 34930 62527 35246 62528
rect 65650 62592 65966 62593
rect 65650 62528 65656 62592
rect 65720 62528 65736 62592
rect 65800 62528 65816 62592
rect 65880 62528 65896 62592
rect 65960 62528 65966 62592
rect 65650 62527 65966 62528
rect 96370 62592 96686 62593
rect 96370 62528 96376 62592
rect 96440 62528 96456 62592
rect 96520 62528 96536 62592
rect 96600 62528 96616 62592
rect 96680 62528 96686 62592
rect 101162 62568 101962 62598
rect 96370 62527 96686 62528
rect 4870 62048 5186 62049
rect 0 61978 800 62008
rect 4870 61984 4876 62048
rect 4940 61984 4956 62048
rect 5020 61984 5036 62048
rect 5100 61984 5116 62048
rect 5180 61984 5186 62048
rect 4870 61983 5186 61984
rect 35590 62048 35906 62049
rect 35590 61984 35596 62048
rect 35660 61984 35676 62048
rect 35740 61984 35756 62048
rect 35820 61984 35836 62048
rect 35900 61984 35906 62048
rect 35590 61983 35906 61984
rect 66310 62048 66626 62049
rect 66310 61984 66316 62048
rect 66380 61984 66396 62048
rect 66460 61984 66476 62048
rect 66540 61984 66556 62048
rect 66620 61984 66626 62048
rect 66310 61983 66626 61984
rect 97030 62048 97346 62049
rect 97030 61984 97036 62048
rect 97100 61984 97116 62048
rect 97180 61984 97196 62048
rect 97260 61984 97276 62048
rect 97340 61984 97346 62048
rect 97030 61983 97346 61984
rect 1485 61978 1551 61981
rect 0 61976 1551 61978
rect 0 61920 1490 61976
rect 1546 61920 1551 61976
rect 0 61918 1551 61920
rect 0 61888 800 61918
rect 1485 61915 1551 61918
rect 100385 61978 100451 61981
rect 101162 61978 101962 62008
rect 100385 61976 101962 61978
rect 100385 61920 100390 61976
rect 100446 61920 101962 61976
rect 100385 61918 101962 61920
rect 100385 61915 100451 61918
rect 101162 61888 101962 61918
rect 4210 61504 4526 61505
rect 4210 61440 4216 61504
rect 4280 61440 4296 61504
rect 4360 61440 4376 61504
rect 4440 61440 4456 61504
rect 4520 61440 4526 61504
rect 4210 61439 4526 61440
rect 34930 61504 35246 61505
rect 34930 61440 34936 61504
rect 35000 61440 35016 61504
rect 35080 61440 35096 61504
rect 35160 61440 35176 61504
rect 35240 61440 35246 61504
rect 34930 61439 35246 61440
rect 65650 61504 65966 61505
rect 65650 61440 65656 61504
rect 65720 61440 65736 61504
rect 65800 61440 65816 61504
rect 65880 61440 65896 61504
rect 65960 61440 65966 61504
rect 65650 61439 65966 61440
rect 96370 61504 96686 61505
rect 96370 61440 96376 61504
rect 96440 61440 96456 61504
rect 96520 61440 96536 61504
rect 96600 61440 96616 61504
rect 96680 61440 96686 61504
rect 96370 61439 96686 61440
rect 841 61434 907 61437
rect 798 61432 907 61434
rect 798 61376 846 61432
rect 902 61376 907 61432
rect 798 61371 907 61376
rect 798 61328 858 61371
rect 0 61238 858 61328
rect 100385 61298 100451 61301
rect 101162 61298 101962 61328
rect 100385 61296 101962 61298
rect 100385 61240 100390 61296
rect 100446 61240 101962 61296
rect 100385 61238 101962 61240
rect 0 61208 800 61238
rect 100385 61235 100451 61238
rect 101162 61208 101962 61238
rect 4870 60960 5186 60961
rect 4870 60896 4876 60960
rect 4940 60896 4956 60960
rect 5020 60896 5036 60960
rect 5100 60896 5116 60960
rect 5180 60896 5186 60960
rect 4870 60895 5186 60896
rect 35590 60960 35906 60961
rect 35590 60896 35596 60960
rect 35660 60896 35676 60960
rect 35740 60896 35756 60960
rect 35820 60896 35836 60960
rect 35900 60896 35906 60960
rect 35590 60895 35906 60896
rect 66310 60960 66626 60961
rect 66310 60896 66316 60960
rect 66380 60896 66396 60960
rect 66460 60896 66476 60960
rect 66540 60896 66556 60960
rect 66620 60896 66626 60960
rect 66310 60895 66626 60896
rect 97030 60960 97346 60961
rect 97030 60896 97036 60960
rect 97100 60896 97116 60960
rect 97180 60896 97196 60960
rect 97260 60896 97276 60960
rect 97340 60896 97346 60960
rect 97030 60895 97346 60896
rect 67582 60692 67588 60756
rect 67652 60754 67658 60756
rect 77109 60754 77175 60757
rect 67652 60752 77175 60754
rect 67652 60696 77114 60752
rect 77170 60696 77175 60752
rect 67652 60694 77175 60696
rect 67652 60692 67658 60694
rect 77109 60691 77175 60694
rect 100385 60618 100451 60621
rect 101162 60618 101962 60648
rect 100385 60616 101962 60618
rect 100385 60560 100390 60616
rect 100446 60560 101962 60616
rect 100385 60558 101962 60560
rect 100385 60555 100451 60558
rect 101162 60528 101962 60558
rect 1302 60416 1458 60417
rect 1302 60352 1308 60416
rect 1372 60352 1388 60416
rect 1452 60352 1458 60416
rect 1302 60351 1458 60352
rect 4210 60416 4526 60417
rect 4210 60352 4216 60416
rect 4280 60352 4296 60416
rect 4360 60352 4376 60416
rect 4440 60352 4456 60416
rect 4520 60352 4526 60416
rect 4210 60351 4526 60352
rect 34930 60416 35246 60417
rect 34930 60352 34936 60416
rect 35000 60352 35016 60416
rect 35080 60352 35096 60416
rect 35160 60352 35176 60416
rect 35240 60352 35246 60416
rect 34930 60351 35246 60352
rect 65650 60416 65966 60417
rect 65650 60352 65656 60416
rect 65720 60352 65736 60416
rect 65800 60352 65816 60416
rect 65880 60352 65896 60416
rect 65960 60352 65966 60416
rect 65650 60351 65966 60352
rect 96370 60416 96686 60417
rect 96370 60352 96376 60416
rect 96440 60352 96456 60416
rect 96520 60352 96536 60416
rect 96600 60352 96616 60416
rect 96680 60352 96686 60416
rect 96370 60351 96686 60352
rect 98926 60416 99242 60417
rect 98926 60352 98932 60416
rect 98996 60352 99012 60416
rect 99076 60352 99092 60416
rect 99156 60352 99172 60416
rect 99236 60352 99242 60416
rect 98926 60351 99242 60352
rect 100385 59938 100451 59941
rect 101162 59938 101962 59968
rect 100385 59936 101962 59938
rect 100385 59880 100390 59936
rect 100446 59880 101962 59936
rect 100385 59878 101962 59880
rect 100385 59875 100451 59878
rect 1670 59872 1826 59873
rect 1670 59808 1676 59872
rect 1740 59808 1756 59872
rect 1820 59808 1826 59872
rect 1670 59807 1826 59808
rect 4870 59872 5186 59873
rect 4870 59808 4876 59872
rect 4940 59808 4956 59872
rect 5020 59808 5036 59872
rect 5100 59808 5116 59872
rect 5180 59808 5186 59872
rect 4870 59807 5186 59808
rect 35590 59872 35906 59873
rect 35590 59808 35596 59872
rect 35660 59808 35676 59872
rect 35740 59808 35756 59872
rect 35820 59808 35836 59872
rect 35900 59808 35906 59872
rect 35590 59807 35906 59808
rect 66310 59872 66626 59873
rect 66310 59808 66316 59872
rect 66380 59808 66396 59872
rect 66460 59808 66476 59872
rect 66540 59808 66556 59872
rect 66620 59808 66626 59872
rect 66310 59807 66626 59808
rect 97030 59872 97346 59873
rect 97030 59808 97036 59872
rect 97100 59808 97116 59872
rect 97180 59808 97196 59872
rect 97260 59808 97276 59872
rect 97340 59808 97346 59872
rect 97030 59807 97346 59808
rect 99662 59872 99978 59873
rect 99662 59808 99668 59872
rect 99732 59808 99748 59872
rect 99812 59808 99828 59872
rect 99892 59808 99908 59872
rect 99972 59808 99978 59872
rect 101162 59848 101962 59878
rect 99662 59807 99978 59808
rect 1302 59328 1458 59329
rect 1302 59264 1308 59328
rect 1372 59264 1388 59328
rect 1452 59264 1458 59328
rect 1302 59263 1458 59264
rect 98926 59328 99242 59329
rect 98926 59264 98932 59328
rect 98996 59264 99012 59328
rect 99076 59264 99092 59328
rect 99156 59264 99172 59328
rect 99236 59264 99242 59328
rect 98926 59263 99242 59264
rect 57462 58788 57468 58852
rect 57532 58850 57538 58852
rect 71773 58850 71839 58853
rect 57532 58848 71839 58850
rect 57532 58792 71778 58848
rect 71834 58792 71839 58848
rect 57532 58790 71839 58792
rect 57532 58788 57538 58790
rect 71773 58787 71839 58790
rect 1670 58784 1826 58785
rect 1670 58720 1676 58784
rect 1740 58720 1756 58784
rect 1820 58720 1826 58784
rect 1670 58719 1826 58720
rect 99662 58784 99978 58785
rect 99662 58720 99668 58784
rect 99732 58720 99748 58784
rect 99812 58720 99828 58784
rect 99892 58720 99908 58784
rect 99972 58720 99978 58784
rect 99662 58719 99978 58720
rect 62614 58652 62620 58716
rect 62684 58714 62690 58716
rect 79501 58714 79567 58717
rect 62684 58712 79567 58714
rect 62684 58656 79506 58712
rect 79562 58656 79567 58712
rect 62684 58654 79567 58656
rect 62684 58652 62690 58654
rect 79501 58651 79567 58654
rect 60038 58516 60044 58580
rect 60108 58578 60114 58580
rect 79133 58578 79199 58581
rect 60108 58576 79199 58578
rect 60108 58520 79138 58576
rect 79194 58520 79199 58576
rect 60108 58518 79199 58520
rect 60108 58516 60114 58518
rect 79133 58515 79199 58518
rect 86125 58578 86191 58581
rect 98269 58578 98335 58581
rect 86125 58576 98335 58578
rect 86125 58520 86130 58576
rect 86186 58520 98274 58576
rect 98330 58520 98335 58576
rect 86125 58518 98335 58520
rect 86125 58515 86191 58518
rect 98269 58515 98335 58518
rect 1302 58240 1458 58241
rect 1302 58176 1308 58240
rect 1372 58176 1388 58240
rect 1452 58176 1458 58240
rect 1302 58175 1458 58176
rect 98926 58240 99242 58241
rect 98926 58176 98932 58240
rect 98996 58176 99012 58240
rect 99076 58176 99092 58240
rect 99156 58176 99172 58240
rect 99236 58176 99242 58240
rect 98926 58175 99242 58176
rect 29177 58170 29243 58173
rect 32565 58170 32571 58172
rect 29177 58168 32571 58170
rect 29177 58112 29182 58168
rect 29238 58112 32571 58168
rect 29177 58110 32571 58112
rect 29177 58107 29243 58110
rect 32565 58108 32571 58110
rect 32635 58108 32641 58172
rect 80136 58108 80142 58172
rect 80206 58170 80212 58172
rect 86125 58170 86191 58173
rect 80206 58168 86191 58170
rect 80206 58112 86130 58168
rect 86186 58112 86191 58168
rect 80206 58110 86191 58112
rect 80206 58108 80212 58110
rect 86125 58107 86191 58110
rect 81304 57972 81310 58036
rect 81374 58034 81380 58036
rect 83917 58034 83983 58037
rect 81374 58032 83983 58034
rect 81374 57976 83922 58032
rect 83978 57976 83983 58032
rect 81374 57974 83983 57976
rect 81374 57972 81380 57974
rect 83917 57971 83983 57974
rect 28165 57898 28231 57901
rect 30069 57898 30075 57900
rect 28165 57896 30075 57898
rect 28165 57840 28170 57896
rect 28226 57840 30075 57896
rect 28165 57838 30075 57840
rect 28165 57835 28231 57838
rect 30069 57836 30075 57838
rect 30139 57836 30145 57900
rect 65013 57836 65019 57900
rect 65083 57898 65089 57900
rect 81801 57898 81867 57901
rect 65083 57896 81867 57898
rect 65083 57840 81806 57896
rect 81862 57840 81867 57896
rect 65083 57838 81867 57840
rect 65083 57836 65089 57838
rect 81801 57835 81867 57838
rect 87873 57898 87939 57901
rect 89852 57898 89858 57900
rect 87873 57896 89858 57898
rect 87873 57840 87878 57896
rect 87934 57840 89858 57896
rect 87873 57838 89858 57840
rect 87873 57835 87939 57838
rect 89852 57836 89858 57838
rect 89922 57898 89928 57900
rect 100109 57898 100175 57901
rect 89922 57896 100175 57898
rect 89922 57840 100114 57896
rect 100170 57840 100175 57896
rect 89922 57838 100175 57840
rect 89922 57836 89928 57838
rect 100109 57835 100175 57838
rect 1670 57696 1826 57697
rect 1670 57632 1676 57696
rect 1740 57632 1756 57696
rect 1820 57632 1826 57696
rect 1670 57631 1826 57632
rect 99662 57696 99978 57697
rect 99662 57632 99668 57696
rect 99732 57632 99748 57696
rect 99812 57632 99828 57696
rect 99892 57632 99908 57696
rect 99972 57632 99978 57696
rect 99662 57631 99978 57632
rect 1302 57152 1458 57153
rect 1302 57088 1308 57152
rect 1372 57088 1388 57152
rect 1452 57088 1458 57152
rect 1302 57087 1458 57088
rect 98926 57152 99242 57153
rect 98926 57088 98932 57152
rect 98996 57088 99012 57152
rect 99076 57088 99092 57152
rect 99156 57088 99172 57152
rect 99236 57088 99242 57152
rect 98926 57087 99242 57088
rect 1670 56608 1826 56609
rect 1670 56544 1676 56608
rect 1740 56544 1756 56608
rect 1820 56544 1826 56608
rect 1670 56543 1826 56544
rect 99662 56608 99978 56609
rect 99662 56544 99668 56608
rect 99732 56544 99748 56608
rect 99812 56544 99828 56608
rect 99892 56544 99908 56608
rect 99972 56544 99978 56608
rect 99662 56543 99978 56544
rect 1302 56064 1458 56065
rect 1302 56000 1308 56064
rect 1372 56000 1388 56064
rect 1452 56000 1458 56064
rect 1302 55999 1458 56000
rect 98926 56064 99242 56065
rect 98926 56000 98932 56064
rect 98996 56000 99012 56064
rect 99076 56000 99092 56064
rect 99156 56000 99172 56064
rect 99236 56000 99242 56064
rect 98926 55999 99242 56000
rect 1670 55520 1826 55521
rect 1670 55456 1676 55520
rect 1740 55456 1756 55520
rect 1820 55456 1826 55520
rect 1670 55455 1826 55456
rect 99662 55520 99978 55521
rect 99662 55456 99668 55520
rect 99732 55456 99748 55520
rect 99812 55456 99828 55520
rect 99892 55456 99908 55520
rect 99972 55456 99978 55520
rect 99662 55455 99978 55456
rect 1302 54976 1458 54977
rect 1302 54912 1308 54976
rect 1372 54912 1388 54976
rect 1452 54912 1458 54976
rect 1302 54911 1458 54912
rect 98926 54976 99242 54977
rect 98926 54912 98932 54976
rect 98996 54912 99012 54976
rect 99076 54912 99092 54976
rect 99156 54912 99172 54976
rect 99236 54912 99242 54976
rect 98926 54911 99242 54912
rect 1670 54432 1826 54433
rect 1670 54368 1676 54432
rect 1740 54368 1756 54432
rect 1820 54368 1826 54432
rect 1670 54367 1826 54368
rect 99662 54432 99978 54433
rect 99662 54368 99668 54432
rect 99732 54368 99748 54432
rect 99812 54368 99828 54432
rect 99892 54368 99908 54432
rect 99972 54368 99978 54432
rect 99662 54367 99978 54368
rect 1302 53888 1458 53889
rect 1302 53824 1308 53888
rect 1372 53824 1388 53888
rect 1452 53824 1458 53888
rect 1302 53823 1458 53824
rect 98926 53888 99242 53889
rect 98926 53824 98932 53888
rect 98996 53824 99012 53888
rect 99076 53824 99092 53888
rect 99156 53824 99172 53888
rect 99236 53824 99242 53888
rect 98926 53823 99242 53824
rect 97073 53818 97139 53821
rect 96478 53816 97139 53818
rect 96478 53768 97078 53816
rect 95956 53760 97078 53768
rect 97134 53760 97139 53816
rect 95956 53758 97139 53760
rect 95956 53708 96538 53758
rect 97073 53755 97139 53758
rect 1670 53344 1826 53345
rect 1670 53280 1676 53344
rect 1740 53280 1756 53344
rect 1820 53280 1826 53344
rect 1670 53279 1826 53280
rect 99662 53344 99978 53345
rect 99662 53280 99668 53344
rect 99732 53280 99748 53344
rect 99812 53280 99828 53344
rect 99892 53280 99908 53344
rect 99972 53280 99978 53344
rect 99662 53279 99978 53280
rect 1302 52800 1458 52801
rect 1302 52736 1308 52800
rect 1372 52736 1388 52800
rect 1452 52736 1458 52800
rect 1302 52735 1458 52736
rect 98926 52800 99242 52801
rect 98926 52736 98932 52800
rect 98996 52736 99012 52800
rect 99076 52736 99092 52800
rect 99156 52736 99172 52800
rect 99236 52736 99242 52800
rect 98926 52735 99242 52736
rect 1670 52256 1826 52257
rect 1670 52192 1676 52256
rect 1740 52192 1756 52256
rect 1820 52192 1826 52256
rect 1670 52191 1826 52192
rect 99662 52256 99978 52257
rect 99662 52192 99668 52256
rect 99732 52192 99748 52256
rect 99812 52192 99828 52256
rect 99892 52192 99908 52256
rect 99972 52192 99978 52256
rect 99662 52191 99978 52192
rect 1302 51712 1458 51713
rect 1302 51648 1308 51712
rect 1372 51648 1388 51712
rect 1452 51648 1458 51712
rect 1302 51647 1458 51648
rect 98926 51712 99242 51713
rect 98926 51648 98932 51712
rect 98996 51648 99012 51712
rect 99076 51648 99092 51712
rect 99156 51648 99172 51712
rect 99236 51648 99242 51712
rect 98926 51647 99242 51648
rect 1670 51168 1826 51169
rect 1670 51104 1676 51168
rect 1740 51104 1756 51168
rect 1820 51104 1826 51168
rect 1670 51103 1826 51104
rect 99662 51168 99978 51169
rect 99662 51104 99668 51168
rect 99732 51104 99748 51168
rect 99812 51104 99828 51168
rect 99892 51104 99908 51168
rect 99972 51104 99978 51168
rect 99662 51103 99978 51104
rect 1302 50624 1458 50625
rect 1302 50560 1308 50624
rect 1372 50560 1388 50624
rect 1452 50560 1458 50624
rect 1302 50559 1458 50560
rect 98926 50624 99242 50625
rect 98926 50560 98932 50624
rect 98996 50560 99012 50624
rect 99076 50560 99092 50624
rect 99156 50560 99172 50624
rect 99236 50560 99242 50624
rect 98926 50559 99242 50560
rect 1670 50080 1826 50081
rect 1670 50016 1676 50080
rect 1740 50016 1756 50080
rect 1820 50016 1826 50080
rect 1670 50015 1826 50016
rect 99662 50080 99978 50081
rect 99662 50016 99668 50080
rect 99732 50016 99748 50080
rect 99812 50016 99828 50080
rect 99892 50016 99908 50080
rect 99972 50016 99978 50080
rect 99662 50015 99978 50016
rect 1302 49536 1458 49537
rect 1302 49472 1308 49536
rect 1372 49472 1388 49536
rect 1452 49472 1458 49536
rect 1302 49471 1458 49472
rect 98926 49536 99242 49537
rect 98926 49472 98932 49536
rect 98996 49472 99012 49536
rect 99076 49472 99092 49536
rect 99156 49472 99172 49536
rect 99236 49472 99242 49536
rect 98926 49471 99242 49472
rect 1670 48992 1826 48993
rect 1670 48928 1676 48992
rect 1740 48928 1756 48992
rect 1820 48928 1826 48992
rect 1670 48927 1826 48928
rect 99662 48992 99978 48993
rect 99662 48928 99668 48992
rect 99732 48928 99748 48992
rect 99812 48928 99828 48992
rect 99892 48928 99908 48992
rect 99972 48928 99978 48992
rect 99662 48927 99978 48928
rect 1302 48448 1458 48449
rect 1302 48384 1308 48448
rect 1372 48384 1388 48448
rect 1452 48384 1458 48448
rect 1302 48383 1458 48384
rect 98926 48448 99242 48449
rect 98926 48384 98932 48448
rect 98996 48384 99012 48448
rect 99076 48384 99092 48448
rect 99156 48384 99172 48448
rect 99236 48384 99242 48448
rect 98926 48383 99242 48384
rect 1670 47904 1826 47905
rect 1670 47840 1676 47904
rect 1740 47840 1756 47904
rect 1820 47840 1826 47904
rect 1670 47839 1826 47840
rect 99662 47904 99978 47905
rect 99662 47840 99668 47904
rect 99732 47840 99748 47904
rect 99812 47840 99828 47904
rect 99892 47840 99908 47904
rect 99972 47840 99978 47904
rect 99662 47839 99978 47840
rect 1302 47360 1458 47361
rect 1302 47296 1308 47360
rect 1372 47296 1388 47360
rect 1452 47296 1458 47360
rect 1302 47295 1458 47296
rect 98926 47360 99242 47361
rect 98926 47296 98932 47360
rect 98996 47296 99012 47360
rect 99076 47296 99092 47360
rect 99156 47296 99172 47360
rect 99236 47296 99242 47360
rect 98926 47295 99242 47296
rect 1670 46816 1826 46817
rect 1670 46752 1676 46816
rect 1740 46752 1756 46816
rect 1820 46752 1826 46816
rect 1670 46751 1826 46752
rect 99662 46816 99978 46817
rect 99662 46752 99668 46816
rect 99732 46752 99748 46816
rect 99812 46752 99828 46816
rect 99892 46752 99908 46816
rect 99972 46752 99978 46816
rect 99662 46751 99978 46752
rect 1302 46272 1458 46273
rect 1302 46208 1308 46272
rect 1372 46208 1388 46272
rect 1452 46208 1458 46272
rect 1302 46207 1458 46208
rect 98926 46272 99242 46273
rect 98926 46208 98932 46272
rect 98996 46208 99012 46272
rect 99076 46208 99092 46272
rect 99156 46208 99172 46272
rect 99236 46208 99242 46272
rect 98926 46207 99242 46208
rect 1670 45728 1826 45729
rect 1670 45664 1676 45728
rect 1740 45664 1756 45728
rect 1820 45664 1826 45728
rect 1670 45663 1826 45664
rect 99662 45728 99978 45729
rect 99662 45664 99668 45728
rect 99732 45664 99748 45728
rect 99812 45664 99828 45728
rect 99892 45664 99908 45728
rect 99972 45664 99978 45728
rect 99662 45663 99978 45664
rect 1302 45184 1458 45185
rect 1302 45120 1308 45184
rect 1372 45120 1388 45184
rect 1452 45120 1458 45184
rect 1302 45119 1458 45120
rect 98926 45184 99242 45185
rect 98926 45120 98932 45184
rect 98996 45120 99012 45184
rect 99076 45120 99092 45184
rect 99156 45120 99172 45184
rect 99236 45120 99242 45184
rect 98926 45119 99242 45120
rect 1670 44640 1826 44641
rect 1670 44576 1676 44640
rect 1740 44576 1756 44640
rect 1820 44576 1826 44640
rect 1670 44575 1826 44576
rect 99662 44640 99978 44641
rect 99662 44576 99668 44640
rect 99732 44576 99748 44640
rect 99812 44576 99828 44640
rect 99892 44576 99908 44640
rect 99972 44576 99978 44640
rect 99662 44575 99978 44576
rect 1302 44096 1458 44097
rect 1302 44032 1308 44096
rect 1372 44032 1388 44096
rect 1452 44032 1458 44096
rect 1302 44031 1458 44032
rect 98926 44096 99242 44097
rect 98926 44032 98932 44096
rect 98996 44032 99012 44096
rect 99076 44032 99092 44096
rect 99156 44032 99172 44096
rect 99236 44032 99242 44096
rect 98926 44031 99242 44032
rect 1670 43552 1826 43553
rect 1670 43488 1676 43552
rect 1740 43488 1756 43552
rect 1820 43488 1826 43552
rect 1670 43487 1826 43488
rect 99662 43552 99978 43553
rect 99662 43488 99668 43552
rect 99732 43488 99748 43552
rect 99812 43488 99828 43552
rect 99892 43488 99908 43552
rect 99972 43488 99978 43552
rect 99662 43487 99978 43488
rect 1302 43008 1458 43009
rect 1302 42944 1308 43008
rect 1372 42944 1388 43008
rect 1452 42944 1458 43008
rect 1302 42943 1458 42944
rect 98926 43008 99242 43009
rect 98926 42944 98932 43008
rect 98996 42944 99012 43008
rect 99076 42944 99092 43008
rect 99156 42944 99172 43008
rect 99236 42944 99242 43008
rect 98926 42943 99242 42944
rect 1670 42464 1826 42465
rect 1670 42400 1676 42464
rect 1740 42400 1756 42464
rect 1820 42400 1826 42464
rect 1670 42399 1826 42400
rect 99662 42464 99978 42465
rect 99662 42400 99668 42464
rect 99732 42400 99748 42464
rect 99812 42400 99828 42464
rect 99892 42400 99908 42464
rect 99972 42400 99978 42464
rect 99662 42399 99978 42400
rect 1302 41920 1458 41921
rect 1302 41856 1308 41920
rect 1372 41856 1388 41920
rect 1452 41856 1458 41920
rect 1302 41855 1458 41856
rect 98926 41920 99242 41921
rect 98926 41856 98932 41920
rect 98996 41856 99012 41920
rect 99076 41856 99092 41920
rect 99156 41856 99172 41920
rect 99236 41856 99242 41920
rect 98926 41855 99242 41856
rect 1670 41376 1826 41377
rect 1670 41312 1676 41376
rect 1740 41312 1756 41376
rect 1820 41312 1826 41376
rect 1670 41311 1826 41312
rect 99662 41376 99978 41377
rect 99662 41312 99668 41376
rect 99732 41312 99748 41376
rect 99812 41312 99828 41376
rect 99892 41312 99908 41376
rect 99972 41312 99978 41376
rect 99662 41311 99978 41312
rect 1302 40832 1458 40833
rect 1302 40768 1308 40832
rect 1372 40768 1388 40832
rect 1452 40768 1458 40832
rect 1302 40767 1458 40768
rect 98926 40832 99242 40833
rect 98926 40768 98932 40832
rect 98996 40768 99012 40832
rect 99076 40768 99092 40832
rect 99156 40768 99172 40832
rect 99236 40768 99242 40832
rect 98926 40767 99242 40768
rect 1670 40288 1826 40289
rect 1670 40224 1676 40288
rect 1740 40224 1756 40288
rect 1820 40224 1826 40288
rect 1670 40223 1826 40224
rect 99662 40288 99978 40289
rect 99662 40224 99668 40288
rect 99732 40224 99748 40288
rect 99812 40224 99828 40288
rect 99892 40224 99908 40288
rect 99972 40224 99978 40288
rect 99662 40223 99978 40224
rect 1302 39744 1458 39745
rect 1302 39680 1308 39744
rect 1372 39680 1388 39744
rect 1452 39680 1458 39744
rect 1302 39679 1458 39680
rect 98926 39744 99242 39745
rect 98926 39680 98932 39744
rect 98996 39680 99012 39744
rect 99076 39680 99092 39744
rect 99156 39680 99172 39744
rect 99236 39680 99242 39744
rect 98926 39679 99242 39680
rect 1670 39200 1826 39201
rect 1670 39136 1676 39200
rect 1740 39136 1756 39200
rect 1820 39136 1826 39200
rect 1670 39135 1826 39136
rect 99662 39200 99978 39201
rect 99662 39136 99668 39200
rect 99732 39136 99748 39200
rect 99812 39136 99828 39200
rect 99892 39136 99908 39200
rect 99972 39136 99978 39200
rect 99662 39135 99978 39136
rect 1302 38656 1458 38657
rect 1302 38592 1308 38656
rect 1372 38592 1388 38656
rect 1452 38592 1458 38656
rect 1302 38591 1458 38592
rect 98926 38656 99242 38657
rect 98926 38592 98932 38656
rect 98996 38592 99012 38656
rect 99076 38592 99092 38656
rect 99156 38592 99172 38656
rect 99236 38592 99242 38656
rect 98926 38591 99242 38592
rect 1670 38112 1826 38113
rect 1670 38048 1676 38112
rect 1740 38048 1756 38112
rect 1820 38048 1826 38112
rect 1670 38047 1826 38048
rect 99662 38112 99978 38113
rect 99662 38048 99668 38112
rect 99732 38048 99748 38112
rect 99812 38048 99828 38112
rect 99892 38048 99908 38112
rect 99972 38048 99978 38112
rect 99662 38047 99978 38048
rect 1302 37568 1458 37569
rect 1302 37504 1308 37568
rect 1372 37504 1388 37568
rect 1452 37504 1458 37568
rect 1302 37503 1458 37504
rect 98926 37568 99242 37569
rect 98926 37504 98932 37568
rect 98996 37504 99012 37568
rect 99076 37504 99092 37568
rect 99156 37504 99172 37568
rect 99236 37504 99242 37568
rect 98926 37503 99242 37504
rect 1670 37024 1826 37025
rect 1670 36960 1676 37024
rect 1740 36960 1756 37024
rect 1820 36960 1826 37024
rect 1670 36959 1826 36960
rect 99662 37024 99978 37025
rect 99662 36960 99668 37024
rect 99732 36960 99748 37024
rect 99812 36960 99828 37024
rect 99892 36960 99908 37024
rect 99972 36960 99978 37024
rect 99662 36959 99978 36960
rect 1302 36480 1458 36481
rect 1302 36416 1308 36480
rect 1372 36416 1388 36480
rect 1452 36416 1458 36480
rect 1302 36415 1458 36416
rect 98926 36480 99242 36481
rect 98926 36416 98932 36480
rect 98996 36416 99012 36480
rect 99076 36416 99092 36480
rect 99156 36416 99172 36480
rect 99236 36416 99242 36480
rect 98926 36415 99242 36416
rect 1670 35936 1826 35937
rect 1670 35872 1676 35936
rect 1740 35872 1756 35936
rect 1820 35872 1826 35936
rect 1670 35871 1826 35872
rect 99662 35936 99978 35937
rect 99662 35872 99668 35936
rect 99732 35872 99748 35936
rect 99812 35872 99828 35936
rect 99892 35872 99908 35936
rect 99972 35872 99978 35936
rect 99662 35871 99978 35872
rect 0 35458 800 35488
rect 0 35398 1226 35458
rect 0 35368 800 35398
rect 1166 35186 1226 35398
rect 1302 35392 1458 35393
rect 1302 35328 1308 35392
rect 1372 35328 1388 35392
rect 1452 35328 1458 35392
rect 1302 35327 1458 35328
rect 98926 35392 99242 35393
rect 98926 35328 98932 35392
rect 98996 35328 99012 35392
rect 99076 35328 99092 35392
rect 99156 35328 99172 35392
rect 99236 35328 99242 35392
rect 98926 35327 99242 35328
rect 3374 35194 4032 35254
rect 3374 35186 3434 35194
rect 1166 35126 3434 35186
rect 1670 34848 1826 34849
rect 1670 34784 1676 34848
rect 1740 34784 1756 34848
rect 1820 34784 1826 34848
rect 1670 34783 1826 34784
rect 99662 34848 99978 34849
rect 99662 34784 99668 34848
rect 99732 34784 99748 34848
rect 99812 34784 99828 34848
rect 99892 34784 99908 34848
rect 99972 34784 99978 34848
rect 99662 34783 99978 34784
rect 1302 34304 1458 34305
rect 1302 34240 1308 34304
rect 1372 34240 1388 34304
rect 1452 34240 1458 34304
rect 1302 34239 1458 34240
rect 98926 34304 99242 34305
rect 98926 34240 98932 34304
rect 98996 34240 99012 34304
rect 99076 34240 99092 34304
rect 99156 34240 99172 34304
rect 99236 34240 99242 34304
rect 98926 34239 99242 34240
rect 1670 33760 1826 33761
rect 1670 33696 1676 33760
rect 1740 33696 1756 33760
rect 1820 33696 1826 33760
rect 1670 33695 1826 33696
rect 99662 33760 99978 33761
rect 99662 33696 99668 33760
rect 99732 33696 99748 33760
rect 99812 33696 99828 33760
rect 99892 33696 99908 33760
rect 99972 33696 99978 33760
rect 99662 33695 99978 33696
rect 2086 33494 4032 33554
rect 0 33418 800 33448
rect 2086 33418 2146 33494
rect 0 33358 2146 33418
rect 0 33328 800 33358
rect 1302 33216 1458 33217
rect 1302 33152 1308 33216
rect 1372 33152 1388 33216
rect 1452 33152 1458 33216
rect 1302 33151 1458 33152
rect 98926 33216 99242 33217
rect 98926 33152 98932 33216
rect 98996 33152 99012 33216
rect 99076 33152 99092 33216
rect 99156 33152 99172 33216
rect 99236 33152 99242 33216
rect 98926 33151 99242 33152
rect 0 32738 800 32768
rect 0 32678 1594 32738
rect 0 32648 800 32678
rect 1534 32466 1594 32678
rect 1670 32672 1826 32673
rect 1670 32608 1676 32672
rect 1740 32608 1756 32672
rect 1820 32608 1826 32672
rect 1670 32607 1826 32608
rect 99662 32672 99978 32673
rect 99662 32608 99668 32672
rect 99732 32608 99748 32672
rect 99812 32608 99828 32672
rect 99892 32608 99908 32672
rect 99972 32608 99978 32672
rect 99662 32607 99978 32608
rect 1534 32426 3434 32466
rect 1534 32406 4032 32426
rect 3374 32366 4032 32406
rect 1302 32128 1458 32129
rect 1302 32064 1308 32128
rect 1372 32064 1388 32128
rect 1452 32064 1458 32128
rect 1302 32063 1458 32064
rect 98926 32128 99242 32129
rect 98926 32064 98932 32128
rect 98996 32064 99012 32128
rect 99076 32064 99092 32128
rect 99156 32064 99172 32128
rect 99236 32064 99242 32128
rect 98926 32063 99242 32064
rect 1670 31584 1826 31585
rect 1670 31520 1676 31584
rect 1740 31520 1756 31584
rect 1820 31520 1826 31584
rect 1670 31519 1826 31520
rect 99662 31584 99978 31585
rect 99662 31520 99668 31584
rect 99732 31520 99748 31584
rect 99812 31520 99828 31584
rect 99892 31520 99908 31584
rect 99972 31520 99978 31584
rect 99662 31519 99978 31520
rect 1302 31040 1458 31041
rect 1302 30976 1308 31040
rect 1372 30976 1388 31040
rect 1452 30976 1458 31040
rect 1302 30975 1458 30976
rect 98926 31040 99242 31041
rect 98926 30976 98932 31040
rect 98996 30976 99012 31040
rect 99076 30976 99092 31040
rect 99156 30976 99172 31040
rect 99236 30976 99242 31040
rect 98926 30975 99242 30976
rect 0 30698 800 30728
rect 3374 30698 4032 30726
rect 0 30666 4032 30698
rect 0 30638 3434 30666
rect 0 30608 800 30638
rect 1670 30496 1826 30497
rect 1670 30432 1676 30496
rect 1740 30432 1756 30496
rect 1820 30432 1826 30496
rect 1670 30431 1826 30432
rect 99662 30496 99978 30497
rect 99662 30432 99668 30496
rect 99732 30432 99748 30496
rect 99812 30432 99828 30496
rect 99892 30432 99908 30496
rect 99972 30432 99978 30496
rect 99662 30431 99978 30432
rect 1302 29952 1458 29953
rect 1302 29888 1308 29952
rect 1372 29888 1388 29952
rect 1452 29888 1458 29952
rect 1302 29887 1458 29888
rect 98926 29952 99242 29953
rect 98926 29888 98932 29952
rect 98996 29888 99012 29952
rect 99076 29888 99092 29952
rect 99156 29888 99172 29952
rect 99236 29888 99242 29952
rect 98926 29887 99242 29888
rect 3374 29610 4032 29643
rect 1534 29583 4032 29610
rect 1534 29550 3434 29583
rect 0 29338 800 29368
rect 1534 29338 1594 29550
rect 1670 29408 1826 29409
rect 1670 29344 1676 29408
rect 1740 29344 1756 29408
rect 1820 29344 1826 29408
rect 1670 29343 1826 29344
rect 99662 29408 99978 29409
rect 99662 29344 99668 29408
rect 99732 29344 99748 29408
rect 99812 29344 99828 29408
rect 99892 29344 99908 29408
rect 99972 29344 99978 29408
rect 99662 29343 99978 29344
rect 0 29278 1594 29338
rect 0 29248 800 29278
rect 1302 28864 1458 28865
rect 1302 28800 1308 28864
rect 1372 28800 1388 28864
rect 1452 28800 1458 28864
rect 1302 28799 1458 28800
rect 98926 28864 99242 28865
rect 98926 28800 98932 28864
rect 98996 28800 99012 28864
rect 99076 28800 99092 28864
rect 99156 28800 99172 28864
rect 99236 28800 99242 28864
rect 98926 28799 99242 28800
rect 1670 28320 1826 28321
rect 1670 28256 1676 28320
rect 1740 28256 1756 28320
rect 1820 28256 1826 28320
rect 1670 28255 1826 28256
rect 99662 28320 99978 28321
rect 99662 28256 99668 28320
rect 99732 28256 99748 28320
rect 99812 28256 99828 28320
rect 99892 28256 99908 28320
rect 99972 28256 99978 28320
rect 99662 28255 99978 28256
rect 0 27978 800 28008
rect 0 27963 3434 27978
rect 0 27918 4032 27963
rect 0 27888 800 27918
rect 3374 27903 4032 27918
rect 1302 27776 1458 27777
rect 1302 27712 1308 27776
rect 1372 27712 1388 27776
rect 1452 27712 1458 27776
rect 1302 27711 1458 27712
rect 98926 27776 99242 27777
rect 98926 27712 98932 27776
rect 98996 27712 99012 27776
rect 99076 27712 99092 27776
rect 99156 27712 99172 27776
rect 99236 27712 99242 27776
rect 98926 27711 99242 27712
rect 1670 27232 1826 27233
rect 1670 27168 1676 27232
rect 1740 27168 1756 27232
rect 1820 27168 1826 27232
rect 1670 27167 1826 27168
rect 99662 27232 99978 27233
rect 99662 27168 99668 27232
rect 99732 27168 99748 27232
rect 99812 27168 99828 27232
rect 99892 27168 99908 27232
rect 99972 27168 99978 27232
rect 99662 27167 99978 27168
rect 1302 26688 1458 26689
rect 1302 26624 1308 26688
rect 1372 26624 1388 26688
rect 1452 26624 1458 26688
rect 1302 26623 1458 26624
rect 98926 26688 99242 26689
rect 98926 26624 98932 26688
rect 98996 26624 99012 26688
rect 99076 26624 99092 26688
rect 99156 26624 99172 26688
rect 99236 26624 99242 26688
rect 98926 26623 99242 26624
rect 1670 26144 1826 26145
rect 1670 26080 1676 26144
rect 1740 26080 1756 26144
rect 1820 26080 1826 26144
rect 1670 26079 1826 26080
rect 99662 26144 99978 26145
rect 99662 26080 99668 26144
rect 99732 26080 99748 26144
rect 99812 26080 99828 26144
rect 99892 26080 99908 26144
rect 99972 26080 99978 26144
rect 99662 26079 99978 26080
rect 100477 25938 100543 25941
rect 101162 25938 101962 25968
rect 100477 25936 101962 25938
rect 100477 25880 100482 25936
rect 100538 25880 101962 25936
rect 100477 25878 101962 25880
rect 100477 25875 100543 25878
rect 101162 25848 101962 25878
rect 1302 25600 1458 25601
rect 1302 25536 1308 25600
rect 1372 25536 1388 25600
rect 1452 25536 1458 25600
rect 1302 25535 1458 25536
rect 98926 25600 99242 25601
rect 98926 25536 98932 25600
rect 98996 25536 99012 25600
rect 99076 25536 99092 25600
rect 99156 25536 99172 25600
rect 99236 25536 99242 25600
rect 98926 25535 99242 25536
rect 1670 25056 1826 25057
rect 1670 24992 1676 25056
rect 1740 24992 1756 25056
rect 1820 24992 1826 25056
rect 1670 24991 1826 24992
rect 99662 25056 99978 25057
rect 99662 24992 99668 25056
rect 99732 24992 99748 25056
rect 99812 24992 99828 25056
rect 99892 24992 99908 25056
rect 99972 24992 99978 25056
rect 99662 24991 99978 24992
rect 1302 24512 1458 24513
rect 1302 24448 1308 24512
rect 1372 24448 1388 24512
rect 1452 24448 1458 24512
rect 1302 24447 1458 24448
rect 98926 24512 99242 24513
rect 98926 24448 98932 24512
rect 98996 24448 99012 24512
rect 99076 24448 99092 24512
rect 99156 24448 99172 24512
rect 99236 24448 99242 24512
rect 98926 24447 99242 24448
rect 1670 23968 1826 23969
rect 1670 23904 1676 23968
rect 1740 23904 1756 23968
rect 1820 23904 1826 23968
rect 1670 23903 1826 23904
rect 99662 23968 99978 23969
rect 99662 23904 99668 23968
rect 99732 23904 99748 23968
rect 99812 23904 99828 23968
rect 99892 23904 99908 23968
rect 99972 23904 99978 23968
rect 99662 23903 99978 23904
rect 1302 23424 1458 23425
rect 1302 23360 1308 23424
rect 1372 23360 1388 23424
rect 1452 23360 1458 23424
rect 1302 23359 1458 23360
rect 98926 23424 99242 23425
rect 98926 23360 98932 23424
rect 98996 23360 99012 23424
rect 99076 23360 99092 23424
rect 99156 23360 99172 23424
rect 99236 23360 99242 23424
rect 98926 23359 99242 23360
rect 1670 22880 1826 22881
rect 1670 22816 1676 22880
rect 1740 22816 1756 22880
rect 1820 22816 1826 22880
rect 1670 22815 1826 22816
rect 99662 22880 99978 22881
rect 99662 22816 99668 22880
rect 99732 22816 99748 22880
rect 99812 22816 99828 22880
rect 99892 22816 99908 22880
rect 99972 22816 99978 22880
rect 99662 22815 99978 22816
rect 1302 22336 1458 22337
rect 1302 22272 1308 22336
rect 1372 22272 1388 22336
rect 1452 22272 1458 22336
rect 1302 22271 1458 22272
rect 98926 22336 99242 22337
rect 98926 22272 98932 22336
rect 98996 22272 99012 22336
rect 99076 22272 99092 22336
rect 99156 22272 99172 22336
rect 99236 22272 99242 22336
rect 98926 22271 99242 22272
rect 1670 21792 1826 21793
rect 1670 21728 1676 21792
rect 1740 21728 1756 21792
rect 1820 21728 1826 21792
rect 1670 21727 1826 21728
rect 99662 21792 99978 21793
rect 99662 21728 99668 21792
rect 99732 21728 99748 21792
rect 99812 21728 99828 21792
rect 99892 21728 99908 21792
rect 99972 21728 99978 21792
rect 99662 21727 99978 21728
rect 1302 21248 1458 21249
rect 1302 21184 1308 21248
rect 1372 21184 1388 21248
rect 1452 21184 1458 21248
rect 1302 21183 1458 21184
rect 98926 21248 99242 21249
rect 98926 21184 98932 21248
rect 98996 21184 99012 21248
rect 99076 21184 99092 21248
rect 99156 21184 99172 21248
rect 99236 21184 99242 21248
rect 98926 21183 99242 21184
rect 1670 20704 1826 20705
rect 1670 20640 1676 20704
rect 1740 20640 1756 20704
rect 1820 20640 1826 20704
rect 1670 20639 1826 20640
rect 99662 20704 99978 20705
rect 99662 20640 99668 20704
rect 99732 20640 99748 20704
rect 99812 20640 99828 20704
rect 99892 20640 99908 20704
rect 99972 20640 99978 20704
rect 99662 20639 99978 20640
rect 1302 20160 1458 20161
rect 1302 20096 1308 20160
rect 1372 20096 1388 20160
rect 1452 20096 1458 20160
rect 1302 20095 1458 20096
rect 98926 20160 99242 20161
rect 98926 20096 98932 20160
rect 98996 20096 99012 20160
rect 99076 20096 99092 20160
rect 99156 20096 99172 20160
rect 99236 20096 99242 20160
rect 98926 20095 99242 20096
rect 1670 19616 1826 19617
rect 1670 19552 1676 19616
rect 1740 19552 1756 19616
rect 1820 19552 1826 19616
rect 1670 19551 1826 19552
rect 99662 19616 99978 19617
rect 99662 19552 99668 19616
rect 99732 19552 99748 19616
rect 99812 19552 99828 19616
rect 99892 19552 99908 19616
rect 99972 19552 99978 19616
rect 99662 19551 99978 19552
rect 98177 19138 98243 19141
rect 96570 19136 98243 19138
rect 96570 19090 98182 19136
rect 95956 19080 98182 19090
rect 98238 19080 98243 19136
rect 95956 19078 98243 19080
rect 1302 19072 1458 19073
rect 1302 19008 1308 19072
rect 1372 19008 1388 19072
rect 1452 19008 1458 19072
rect 95956 19030 96630 19078
rect 98177 19075 98243 19078
rect 98926 19072 99242 19073
rect 1302 19007 1458 19008
rect 98926 19008 98932 19072
rect 98996 19008 99012 19072
rect 99076 19008 99092 19072
rect 99156 19008 99172 19072
rect 99236 19008 99242 19072
rect 98926 19007 99242 19008
rect 1670 18528 1826 18529
rect 1670 18464 1676 18528
rect 1740 18464 1756 18528
rect 1820 18464 1826 18528
rect 1670 18463 1826 18464
rect 99662 18528 99978 18529
rect 99662 18464 99668 18528
rect 99732 18464 99748 18528
rect 99812 18464 99828 18528
rect 99892 18464 99908 18528
rect 99972 18464 99978 18528
rect 99662 18463 99978 18464
rect 1302 17984 1458 17985
rect 1302 17920 1308 17984
rect 1372 17920 1388 17984
rect 1452 17920 1458 17984
rect 1302 17919 1458 17920
rect 98926 17984 99242 17985
rect 98926 17920 98932 17984
rect 98996 17920 99012 17984
rect 99076 17920 99092 17984
rect 99156 17920 99172 17984
rect 99236 17920 99242 17984
rect 98926 17919 99242 17920
rect 1670 17440 1826 17441
rect 1670 17376 1676 17440
rect 1740 17376 1756 17440
rect 1820 17376 1826 17440
rect 99662 17440 99978 17441
rect 1670 17375 1826 17376
rect 95956 17370 96630 17390
rect 99662 17376 99668 17440
rect 99732 17376 99748 17440
rect 99812 17376 99828 17440
rect 99892 17376 99908 17440
rect 99972 17376 99978 17440
rect 99662 17375 99978 17376
rect 99373 17370 99439 17373
rect 95956 17368 99439 17370
rect 95956 17330 99378 17368
rect 96570 17312 99378 17330
rect 99434 17312 99439 17368
rect 96570 17310 99439 17312
rect 99373 17307 99439 17310
rect 1302 16896 1458 16897
rect 1302 16832 1308 16896
rect 1372 16832 1388 16896
rect 1452 16832 1458 16896
rect 1302 16831 1458 16832
rect 98926 16896 99242 16897
rect 98926 16832 98932 16896
rect 98996 16832 99012 16896
rect 99076 16832 99092 16896
rect 99156 16832 99172 16896
rect 99236 16832 99242 16896
rect 98926 16831 99242 16832
rect 1670 16352 1826 16353
rect 1670 16288 1676 16352
rect 1740 16288 1756 16352
rect 1820 16288 1826 16352
rect 1670 16287 1826 16288
rect 99662 16352 99978 16353
rect 99662 16288 99668 16352
rect 99732 16288 99748 16352
rect 99812 16288 99828 16352
rect 99892 16288 99908 16352
rect 99972 16288 99978 16352
rect 99662 16287 99978 16288
rect 98545 16282 98611 16285
rect 96478 16280 98611 16282
rect 96478 16262 98550 16280
rect 95956 16224 98550 16262
rect 98606 16224 98611 16280
rect 95956 16222 98611 16224
rect 95956 16202 96538 16222
rect 98545 16219 98611 16222
rect 1302 15808 1458 15809
rect 1302 15744 1308 15808
rect 1372 15744 1388 15808
rect 1452 15744 1458 15808
rect 1302 15743 1458 15744
rect 98926 15808 99242 15809
rect 98926 15744 98932 15808
rect 98996 15744 99012 15808
rect 99076 15744 99092 15808
rect 99156 15744 99172 15808
rect 99236 15744 99242 15808
rect 98926 15743 99242 15744
rect 1670 15264 1826 15265
rect 1670 15200 1676 15264
rect 1740 15200 1756 15264
rect 1820 15200 1826 15264
rect 1670 15199 1826 15200
rect 99662 15264 99978 15265
rect 99662 15200 99668 15264
rect 99732 15200 99748 15264
rect 99812 15200 99828 15264
rect 99892 15200 99908 15264
rect 99972 15200 99978 15264
rect 99662 15199 99978 15200
rect 1302 14720 1458 14721
rect 1302 14656 1308 14720
rect 1372 14656 1388 14720
rect 1452 14656 1458 14720
rect 1302 14655 1458 14656
rect 98926 14720 99242 14721
rect 98926 14656 98932 14720
rect 98996 14656 99012 14720
rect 99076 14656 99092 14720
rect 99156 14656 99172 14720
rect 99236 14656 99242 14720
rect 98926 14655 99242 14656
rect 1670 14176 1826 14177
rect 1670 14112 1676 14176
rect 1740 14112 1756 14176
rect 1820 14112 1826 14176
rect 1670 14111 1826 14112
rect 99662 14176 99978 14177
rect 99662 14112 99668 14176
rect 99732 14112 99748 14176
rect 99812 14112 99828 14176
rect 99892 14112 99908 14176
rect 99972 14112 99978 14176
rect 99662 14111 99978 14112
rect 1302 13632 1458 13633
rect 1302 13568 1308 13632
rect 1372 13568 1388 13632
rect 1452 13568 1458 13632
rect 1302 13567 1458 13568
rect 98926 13632 99242 13633
rect 98926 13568 98932 13632
rect 98996 13568 99012 13632
rect 99076 13568 99092 13632
rect 99156 13568 99172 13632
rect 99236 13568 99242 13632
rect 98926 13567 99242 13568
rect 1670 13088 1826 13089
rect 1670 13024 1676 13088
rect 1740 13024 1756 13088
rect 1820 13024 1826 13088
rect 1670 13023 1826 13024
rect 99662 13088 99978 13089
rect 99662 13024 99668 13088
rect 99732 13024 99748 13088
rect 99812 13024 99828 13088
rect 99892 13024 99908 13088
rect 99972 13024 99978 13088
rect 99662 13023 99978 13024
rect 1302 12544 1458 12545
rect 1302 12480 1308 12544
rect 1372 12480 1388 12544
rect 1452 12480 1458 12544
rect 1302 12479 1458 12480
rect 98926 12544 99242 12545
rect 98926 12480 98932 12544
rect 98996 12480 99012 12544
rect 99076 12480 99092 12544
rect 99156 12480 99172 12544
rect 99236 12480 99242 12544
rect 98926 12479 99242 12480
rect 1670 12000 1826 12001
rect 1670 11936 1676 12000
rect 1740 11936 1756 12000
rect 1820 11936 1826 12000
rect 1670 11935 1826 11936
rect 99662 12000 99978 12001
rect 99662 11936 99668 12000
rect 99732 11936 99748 12000
rect 99812 11936 99828 12000
rect 99892 11936 99908 12000
rect 99972 11936 99978 12000
rect 99662 11935 99978 11936
rect 1302 11456 1458 11457
rect 1302 11392 1308 11456
rect 1372 11392 1388 11456
rect 1452 11392 1458 11456
rect 1302 11391 1458 11392
rect 98926 11456 99242 11457
rect 98926 11392 98932 11456
rect 98996 11392 99012 11456
rect 99076 11392 99092 11456
rect 99156 11392 99172 11456
rect 99236 11392 99242 11456
rect 98926 11391 99242 11392
rect 1670 10912 1826 10913
rect 1670 10848 1676 10912
rect 1740 10848 1756 10912
rect 1820 10848 1826 10912
rect 1670 10847 1826 10848
rect 99662 10912 99978 10913
rect 99662 10848 99668 10912
rect 99732 10848 99748 10912
rect 99812 10848 99828 10912
rect 99892 10848 99908 10912
rect 99972 10848 99978 10912
rect 99662 10847 99978 10848
rect 1302 10368 1458 10369
rect 1302 10304 1308 10368
rect 1372 10304 1388 10368
rect 1452 10304 1458 10368
rect 1302 10303 1458 10304
rect 98926 10368 99242 10369
rect 98926 10304 98932 10368
rect 98996 10304 99012 10368
rect 99076 10304 99092 10368
rect 99156 10304 99172 10368
rect 99236 10304 99242 10368
rect 98926 10303 99242 10304
rect 1670 9824 1826 9825
rect 1670 9760 1676 9824
rect 1740 9760 1756 9824
rect 1820 9760 1826 9824
rect 1670 9759 1826 9760
rect 99662 9824 99978 9825
rect 99662 9760 99668 9824
rect 99732 9760 99748 9824
rect 99812 9760 99828 9824
rect 99892 9760 99908 9824
rect 99972 9760 99978 9824
rect 99662 9759 99978 9760
rect 0 9618 800 9648
rect 0 9558 3434 9618
rect 0 9528 800 9558
rect 3374 9483 3434 9558
rect 3374 9423 4032 9483
rect 1302 9280 1458 9281
rect 1302 9216 1308 9280
rect 1372 9216 1388 9280
rect 1452 9216 1458 9280
rect 1302 9215 1458 9216
rect 98926 9280 99242 9281
rect 98926 9216 98932 9280
rect 98996 9216 99012 9280
rect 99076 9216 99092 9280
rect 99156 9216 99172 9280
rect 99236 9216 99242 9280
rect 98926 9215 99242 9216
rect 1670 8736 1826 8737
rect 1670 8672 1676 8736
rect 1740 8672 1756 8736
rect 1820 8672 1826 8736
rect 1670 8671 1826 8672
rect 99662 8736 99978 8737
rect 99662 8672 99668 8736
rect 99732 8672 99748 8736
rect 99812 8672 99828 8736
rect 99892 8672 99908 8736
rect 99972 8672 99978 8736
rect 99662 8671 99978 8672
rect 1302 8192 1458 8193
rect 1302 8128 1308 8192
rect 1372 8128 1388 8192
rect 1452 8128 1458 8192
rect 1302 8127 1458 8128
rect 98926 8192 99242 8193
rect 98926 8128 98932 8192
rect 98996 8128 99012 8192
rect 99076 8128 99092 8192
rect 99156 8128 99172 8192
rect 99236 8128 99242 8192
rect 98926 8127 99242 8128
rect 1670 7648 1826 7649
rect 1670 7584 1676 7648
rect 1740 7584 1756 7648
rect 1820 7584 1826 7648
rect 1670 7583 1826 7584
rect 99662 7648 99978 7649
rect 99662 7584 99668 7648
rect 99732 7584 99748 7648
rect 99812 7584 99828 7648
rect 99892 7584 99908 7648
rect 99972 7584 99978 7648
rect 99662 7583 99978 7584
rect 1302 7104 1458 7105
rect 1302 7040 1308 7104
rect 1372 7040 1388 7104
rect 1452 7040 1458 7104
rect 1302 7039 1458 7040
rect 98926 7104 99242 7105
rect 98926 7040 98932 7104
rect 98996 7040 99012 7104
rect 99076 7040 99092 7104
rect 99156 7040 99172 7104
rect 99236 7040 99242 7104
rect 98926 7039 99242 7040
rect 1670 6560 1826 6561
rect 1670 6496 1676 6560
rect 1740 6496 1756 6560
rect 1820 6496 1826 6560
rect 1670 6495 1826 6496
rect 99662 6560 99978 6561
rect 99662 6496 99668 6560
rect 99732 6496 99748 6560
rect 99812 6496 99828 6560
rect 99892 6496 99908 6560
rect 99972 6496 99978 6560
rect 99662 6495 99978 6496
rect 1302 6016 1458 6017
rect 1302 5952 1308 6016
rect 1372 5952 1388 6016
rect 1452 5952 1458 6016
rect 1302 5951 1458 5952
rect 98926 6016 99242 6017
rect 98926 5952 98932 6016
rect 98996 5952 99012 6016
rect 99076 5952 99092 6016
rect 99156 5952 99172 6016
rect 99236 5952 99242 6016
rect 98926 5951 99242 5952
rect 1670 5472 1826 5473
rect 1670 5408 1676 5472
rect 1740 5408 1756 5472
rect 1820 5408 1826 5472
rect 1670 5407 1826 5408
rect 99662 5472 99978 5473
rect 99662 5408 99668 5472
rect 99732 5408 99748 5472
rect 99812 5408 99828 5472
rect 99892 5408 99908 5472
rect 99972 5408 99978 5472
rect 99662 5407 99978 5408
rect 1302 4928 1458 4929
rect 1302 4864 1308 4928
rect 1372 4864 1388 4928
rect 1452 4864 1458 4928
rect 1302 4863 1458 4864
rect 98926 4928 99242 4929
rect 98926 4864 98932 4928
rect 98996 4864 99012 4928
rect 99076 4864 99092 4928
rect 99156 4864 99172 4928
rect 99236 4864 99242 4928
rect 98926 4863 99242 4864
rect 1670 4384 1826 4385
rect 1670 4320 1676 4384
rect 1740 4320 1756 4384
rect 1820 4320 1826 4384
rect 1670 4319 1826 4320
rect 99662 4384 99978 4385
rect 99662 4320 99668 4384
rect 99732 4320 99748 4384
rect 99812 4320 99828 4384
rect 99892 4320 99908 4384
rect 99972 4320 99978 4384
rect 99662 4319 99978 4320
rect 97257 4178 97323 4181
rect 101162 4178 101962 4208
rect 97257 4176 101962 4178
rect 97257 4120 97262 4176
rect 97318 4120 101962 4176
rect 97257 4118 101962 4120
rect 97257 4115 97323 4118
rect 101162 4088 101962 4118
rect 2681 3906 2747 3909
rect 10052 3906 10058 3908
rect 2681 3904 10058 3906
rect 2681 3848 2686 3904
rect 2742 3848 10058 3904
rect 2681 3846 10058 3848
rect 2681 3843 2747 3846
rect 10052 3844 10058 3846
rect 10122 3844 10128 3908
rect 84808 3844 84814 3908
rect 84878 3906 84884 3908
rect 97993 3906 98059 3909
rect 84878 3904 98059 3906
rect 84878 3848 97998 3904
rect 98054 3848 98059 3904
rect 84878 3846 98059 3848
rect 84878 3844 84884 3846
rect 97993 3843 98059 3846
rect 1302 3840 1458 3841
rect 1302 3776 1308 3840
rect 1372 3776 1388 3840
rect 1452 3776 1458 3840
rect 1302 3775 1458 3776
rect 98926 3840 99242 3841
rect 98926 3776 98932 3840
rect 98996 3776 99012 3840
rect 99076 3776 99092 3840
rect 99156 3776 99172 3840
rect 99236 3776 99242 3840
rect 98926 3775 99242 3776
rect 84659 3708 84665 3772
rect 84729 3770 84735 3772
rect 97533 3770 97599 3773
rect 84729 3768 97599 3770
rect 84729 3712 97538 3768
rect 97594 3712 97599 3768
rect 84729 3710 97599 3712
rect 84729 3708 84735 3710
rect 97533 3707 97599 3710
rect 84521 3572 84527 3636
rect 84591 3634 84597 3636
rect 97349 3634 97415 3637
rect 84591 3632 97415 3634
rect 84591 3576 97354 3632
rect 97410 3576 97415 3632
rect 84591 3574 97415 3576
rect 84591 3572 84597 3574
rect 97349 3571 97415 3574
rect 17401 3500 17467 3501
rect 17401 3496 17438 3500
rect 17502 3498 17508 3500
rect 17401 3440 17406 3496
rect 17401 3436 17438 3440
rect 17502 3438 17558 3498
rect 17502 3436 17508 3438
rect 19768 3436 19774 3500
rect 19838 3498 19844 3500
rect 19977 3498 20043 3501
rect 19838 3496 20043 3498
rect 19838 3440 19982 3496
rect 20038 3440 20043 3496
rect 19838 3438 20043 3440
rect 19838 3436 19844 3438
rect 17401 3435 17467 3436
rect 19977 3435 20043 3438
rect 20621 3498 20687 3501
rect 20936 3498 20942 3500
rect 20621 3496 20942 3498
rect 20621 3440 20626 3496
rect 20682 3440 20942 3496
rect 20621 3438 20942 3440
rect 20621 3435 20687 3438
rect 20936 3436 20942 3438
rect 21006 3436 21012 3500
rect 21909 3498 21975 3501
rect 24485 3500 24551 3501
rect 22104 3498 22110 3500
rect 21909 3496 22110 3498
rect 21909 3440 21914 3496
rect 21970 3440 22110 3496
rect 21909 3438 22110 3440
rect 21909 3435 21975 3438
rect 22104 3436 22110 3438
rect 22174 3436 22180 3500
rect 24440 3498 24446 3500
rect 24394 3438 24446 3498
rect 24510 3496 24551 3500
rect 24546 3440 24551 3496
rect 24440 3436 24446 3438
rect 24510 3436 24551 3440
rect 25608 3436 25614 3500
rect 25678 3498 25684 3500
rect 25773 3498 25839 3501
rect 25678 3496 25839 3498
rect 25678 3440 25778 3496
rect 25834 3440 25839 3496
rect 25678 3438 25839 3440
rect 25678 3436 25684 3438
rect 24485 3435 24551 3436
rect 25773 3435 25839 3438
rect 26776 3436 26782 3500
rect 26846 3498 26852 3500
rect 27061 3498 27127 3501
rect 26846 3496 27127 3498
rect 26846 3440 27066 3496
rect 27122 3440 27127 3496
rect 26846 3438 27127 3440
rect 26846 3436 26852 3438
rect 27061 3435 27127 3438
rect 27705 3498 27771 3501
rect 30281 3500 30347 3501
rect 27930 3498 27936 3500
rect 27705 3496 27936 3498
rect 27705 3440 27710 3496
rect 27766 3440 27936 3496
rect 27705 3438 27936 3440
rect 27705 3435 27771 3438
rect 27930 3436 27936 3438
rect 28000 3436 28006 3500
rect 30280 3436 30286 3500
rect 30350 3498 30356 3500
rect 33501 3498 33567 3501
rect 33784 3498 33790 3500
rect 30350 3438 30438 3498
rect 33501 3496 33790 3498
rect 33501 3440 33506 3496
rect 33562 3440 33790 3496
rect 33501 3438 33790 3440
rect 30350 3436 30356 3438
rect 30281 3435 30347 3436
rect 33501 3435 33567 3438
rect 33784 3436 33790 3438
rect 33854 3436 33860 3500
rect 34789 3498 34855 3501
rect 34952 3498 34958 3500
rect 34789 3496 34958 3498
rect 34789 3440 34794 3496
rect 34850 3440 34958 3496
rect 34789 3438 34958 3440
rect 34789 3435 34855 3438
rect 34952 3436 34958 3438
rect 35022 3436 35028 3500
rect 1670 3296 1826 3297
rect 1670 3232 1676 3296
rect 1740 3232 1756 3296
rect 1820 3232 1826 3296
rect 1670 3231 1826 3232
rect 99662 3296 99978 3297
rect 99662 3232 99668 3296
rect 99732 3232 99748 3296
rect 99812 3232 99828 3296
rect 99892 3232 99908 3296
rect 99972 3232 99978 3296
rect 99662 3231 99978 3232
rect 18689 2820 18755 2821
rect 18638 2818 18644 2820
rect 18598 2758 18644 2818
rect 18708 2816 18755 2820
rect 18750 2760 18755 2816
rect 18638 2756 18644 2758
rect 18708 2756 18755 2760
rect 18689 2755 18755 2756
rect 23197 2820 23263 2821
rect 23197 2816 23244 2820
rect 23308 2818 23314 2820
rect 28993 2818 29059 2821
rect 31569 2820 31635 2821
rect 29126 2818 29132 2820
rect 23197 2760 23202 2816
rect 23197 2756 23244 2760
rect 23308 2758 23354 2818
rect 28993 2816 29132 2818
rect 28993 2760 28998 2816
rect 29054 2760 29132 2816
rect 28993 2758 29132 2760
rect 23308 2756 23314 2758
rect 23197 2755 23263 2756
rect 28993 2755 29059 2758
rect 29126 2756 29132 2758
rect 29196 2756 29202 2820
rect 31518 2818 31524 2820
rect 31478 2758 31524 2818
rect 31588 2816 31635 2820
rect 31630 2760 31635 2816
rect 31518 2756 31524 2758
rect 31588 2756 31635 2760
rect 32622 2756 32628 2820
rect 32692 2818 32698 2820
rect 32857 2818 32923 2821
rect 36077 2820 36143 2821
rect 36077 2818 36124 2820
rect 32692 2816 32923 2818
rect 32692 2760 32862 2816
rect 32918 2760 32923 2816
rect 32692 2758 32923 2760
rect 36032 2816 36124 2818
rect 36032 2760 36082 2816
rect 36032 2758 36124 2760
rect 32692 2756 32698 2758
rect 31569 2755 31635 2756
rect 32857 2755 32923 2758
rect 36077 2756 36124 2758
rect 36188 2756 36194 2820
rect 37222 2756 37228 2820
rect 37292 2818 37298 2820
rect 37365 2818 37431 2821
rect 37292 2816 37431 2818
rect 37292 2760 37370 2816
rect 37426 2760 37431 2816
rect 37292 2758 37431 2760
rect 37292 2756 37298 2758
rect 36077 2755 36143 2756
rect 37365 2755 37431 2758
rect 1302 2752 1458 2753
rect 1302 2688 1308 2752
rect 1372 2688 1388 2752
rect 1452 2688 1458 2752
rect 1302 2687 1458 2688
rect 98926 2752 99242 2753
rect 98926 2688 98932 2752
rect 98996 2688 99012 2752
rect 99076 2688 99092 2752
rect 99156 2688 99172 2752
rect 99236 2688 99242 2752
rect 98926 2687 99242 2688
rect 1670 2208 1826 2209
rect 1670 2144 1676 2208
rect 1740 2144 1756 2208
rect 1820 2144 1826 2208
rect 1670 2143 1826 2144
rect 99662 2208 99978 2209
rect 99662 2144 99668 2208
rect 99732 2144 99748 2208
rect 99812 2144 99828 2208
rect 99892 2144 99908 2208
rect 99972 2144 99978 2208
rect 99662 2143 99978 2144
<< via3 >>
rect 4216 101756 4280 101760
rect 4216 101700 4220 101756
rect 4220 101700 4276 101756
rect 4276 101700 4280 101756
rect 4216 101696 4280 101700
rect 4296 101756 4360 101760
rect 4296 101700 4300 101756
rect 4300 101700 4356 101756
rect 4356 101700 4360 101756
rect 4296 101696 4360 101700
rect 4376 101756 4440 101760
rect 4376 101700 4380 101756
rect 4380 101700 4436 101756
rect 4436 101700 4440 101756
rect 4376 101696 4440 101700
rect 4456 101756 4520 101760
rect 4456 101700 4460 101756
rect 4460 101700 4516 101756
rect 4516 101700 4520 101756
rect 4456 101696 4520 101700
rect 34936 101756 35000 101760
rect 34936 101700 34940 101756
rect 34940 101700 34996 101756
rect 34996 101700 35000 101756
rect 34936 101696 35000 101700
rect 35016 101756 35080 101760
rect 35016 101700 35020 101756
rect 35020 101700 35076 101756
rect 35076 101700 35080 101756
rect 35016 101696 35080 101700
rect 35096 101756 35160 101760
rect 35096 101700 35100 101756
rect 35100 101700 35156 101756
rect 35156 101700 35160 101756
rect 35096 101696 35160 101700
rect 35176 101756 35240 101760
rect 35176 101700 35180 101756
rect 35180 101700 35236 101756
rect 35236 101700 35240 101756
rect 35176 101696 35240 101700
rect 65656 101756 65720 101760
rect 65656 101700 65660 101756
rect 65660 101700 65716 101756
rect 65716 101700 65720 101756
rect 65656 101696 65720 101700
rect 65736 101756 65800 101760
rect 65736 101700 65740 101756
rect 65740 101700 65796 101756
rect 65796 101700 65800 101756
rect 65736 101696 65800 101700
rect 65816 101756 65880 101760
rect 65816 101700 65820 101756
rect 65820 101700 65876 101756
rect 65876 101700 65880 101756
rect 65816 101696 65880 101700
rect 65896 101756 65960 101760
rect 65896 101700 65900 101756
rect 65900 101700 65956 101756
rect 65956 101700 65960 101756
rect 65896 101696 65960 101700
rect 96376 101756 96440 101760
rect 96376 101700 96380 101756
rect 96380 101700 96436 101756
rect 96436 101700 96440 101756
rect 96376 101696 96440 101700
rect 96456 101756 96520 101760
rect 96456 101700 96460 101756
rect 96460 101700 96516 101756
rect 96516 101700 96520 101756
rect 96456 101696 96520 101700
rect 96536 101756 96600 101760
rect 96536 101700 96540 101756
rect 96540 101700 96596 101756
rect 96596 101700 96600 101756
rect 96536 101696 96600 101700
rect 96616 101756 96680 101760
rect 96616 101700 96620 101756
rect 96620 101700 96676 101756
rect 96676 101700 96680 101756
rect 96616 101696 96680 101700
rect 4876 101212 4940 101216
rect 4876 101156 4880 101212
rect 4880 101156 4936 101212
rect 4936 101156 4940 101212
rect 4876 101152 4940 101156
rect 4956 101212 5020 101216
rect 4956 101156 4960 101212
rect 4960 101156 5016 101212
rect 5016 101156 5020 101212
rect 4956 101152 5020 101156
rect 5036 101212 5100 101216
rect 5036 101156 5040 101212
rect 5040 101156 5096 101212
rect 5096 101156 5100 101212
rect 5036 101152 5100 101156
rect 5116 101212 5180 101216
rect 5116 101156 5120 101212
rect 5120 101156 5176 101212
rect 5176 101156 5180 101212
rect 5116 101152 5180 101156
rect 35596 101212 35660 101216
rect 35596 101156 35600 101212
rect 35600 101156 35656 101212
rect 35656 101156 35660 101212
rect 35596 101152 35660 101156
rect 35676 101212 35740 101216
rect 35676 101156 35680 101212
rect 35680 101156 35736 101212
rect 35736 101156 35740 101212
rect 35676 101152 35740 101156
rect 35756 101212 35820 101216
rect 35756 101156 35760 101212
rect 35760 101156 35816 101212
rect 35816 101156 35820 101212
rect 35756 101152 35820 101156
rect 35836 101212 35900 101216
rect 35836 101156 35840 101212
rect 35840 101156 35896 101212
rect 35896 101156 35900 101212
rect 35836 101152 35900 101156
rect 66316 101212 66380 101216
rect 66316 101156 66320 101212
rect 66320 101156 66376 101212
rect 66376 101156 66380 101212
rect 66316 101152 66380 101156
rect 66396 101212 66460 101216
rect 66396 101156 66400 101212
rect 66400 101156 66456 101212
rect 66456 101156 66460 101212
rect 66396 101152 66460 101156
rect 66476 101212 66540 101216
rect 66476 101156 66480 101212
rect 66480 101156 66536 101212
rect 66536 101156 66540 101212
rect 66476 101152 66540 101156
rect 66556 101212 66620 101216
rect 66556 101156 66560 101212
rect 66560 101156 66616 101212
rect 66616 101156 66620 101212
rect 66556 101152 66620 101156
rect 97036 101212 97100 101216
rect 97036 101156 97040 101212
rect 97040 101156 97096 101212
rect 97096 101156 97100 101212
rect 97036 101152 97100 101156
rect 97116 101212 97180 101216
rect 97116 101156 97120 101212
rect 97120 101156 97176 101212
rect 97176 101156 97180 101212
rect 97116 101152 97180 101156
rect 97196 101212 97260 101216
rect 97196 101156 97200 101212
rect 97200 101156 97256 101212
rect 97256 101156 97260 101212
rect 97196 101152 97260 101156
rect 97276 101212 97340 101216
rect 97276 101156 97280 101212
rect 97280 101156 97336 101212
rect 97336 101156 97340 101212
rect 97276 101152 97340 101156
rect 4216 100668 4280 100672
rect 4216 100612 4220 100668
rect 4220 100612 4276 100668
rect 4276 100612 4280 100668
rect 4216 100608 4280 100612
rect 4296 100668 4360 100672
rect 4296 100612 4300 100668
rect 4300 100612 4356 100668
rect 4356 100612 4360 100668
rect 4296 100608 4360 100612
rect 4376 100668 4440 100672
rect 4376 100612 4380 100668
rect 4380 100612 4436 100668
rect 4436 100612 4440 100668
rect 4376 100608 4440 100612
rect 4456 100668 4520 100672
rect 4456 100612 4460 100668
rect 4460 100612 4516 100668
rect 4516 100612 4520 100668
rect 4456 100608 4520 100612
rect 34936 100668 35000 100672
rect 34936 100612 34940 100668
rect 34940 100612 34996 100668
rect 34996 100612 35000 100668
rect 34936 100608 35000 100612
rect 35016 100668 35080 100672
rect 35016 100612 35020 100668
rect 35020 100612 35076 100668
rect 35076 100612 35080 100668
rect 35016 100608 35080 100612
rect 35096 100668 35160 100672
rect 35096 100612 35100 100668
rect 35100 100612 35156 100668
rect 35156 100612 35160 100668
rect 35096 100608 35160 100612
rect 35176 100668 35240 100672
rect 35176 100612 35180 100668
rect 35180 100612 35236 100668
rect 35236 100612 35240 100668
rect 35176 100608 35240 100612
rect 65656 100668 65720 100672
rect 65656 100612 65660 100668
rect 65660 100612 65716 100668
rect 65716 100612 65720 100668
rect 65656 100608 65720 100612
rect 65736 100668 65800 100672
rect 65736 100612 65740 100668
rect 65740 100612 65796 100668
rect 65796 100612 65800 100668
rect 65736 100608 65800 100612
rect 65816 100668 65880 100672
rect 65816 100612 65820 100668
rect 65820 100612 65876 100668
rect 65876 100612 65880 100668
rect 65816 100608 65880 100612
rect 65896 100668 65960 100672
rect 65896 100612 65900 100668
rect 65900 100612 65956 100668
rect 65956 100612 65960 100668
rect 65896 100608 65960 100612
rect 96376 100668 96440 100672
rect 96376 100612 96380 100668
rect 96380 100612 96436 100668
rect 96436 100612 96440 100668
rect 96376 100608 96440 100612
rect 96456 100668 96520 100672
rect 96456 100612 96460 100668
rect 96460 100612 96516 100668
rect 96516 100612 96520 100668
rect 96456 100608 96520 100612
rect 96536 100668 96600 100672
rect 96536 100612 96540 100668
rect 96540 100612 96596 100668
rect 96596 100612 96600 100668
rect 96536 100608 96600 100612
rect 96616 100668 96680 100672
rect 96616 100612 96620 100668
rect 96620 100612 96676 100668
rect 96676 100612 96680 100668
rect 96616 100608 96680 100612
rect 4876 100124 4940 100128
rect 4876 100068 4880 100124
rect 4880 100068 4936 100124
rect 4936 100068 4940 100124
rect 4876 100064 4940 100068
rect 4956 100124 5020 100128
rect 4956 100068 4960 100124
rect 4960 100068 5016 100124
rect 5016 100068 5020 100124
rect 4956 100064 5020 100068
rect 5036 100124 5100 100128
rect 5036 100068 5040 100124
rect 5040 100068 5096 100124
rect 5096 100068 5100 100124
rect 5036 100064 5100 100068
rect 5116 100124 5180 100128
rect 5116 100068 5120 100124
rect 5120 100068 5176 100124
rect 5176 100068 5180 100124
rect 5116 100064 5180 100068
rect 35596 100124 35660 100128
rect 35596 100068 35600 100124
rect 35600 100068 35656 100124
rect 35656 100068 35660 100124
rect 35596 100064 35660 100068
rect 35676 100124 35740 100128
rect 35676 100068 35680 100124
rect 35680 100068 35736 100124
rect 35736 100068 35740 100124
rect 35676 100064 35740 100068
rect 35756 100124 35820 100128
rect 35756 100068 35760 100124
rect 35760 100068 35816 100124
rect 35816 100068 35820 100124
rect 35756 100064 35820 100068
rect 35836 100124 35900 100128
rect 35836 100068 35840 100124
rect 35840 100068 35896 100124
rect 35896 100068 35900 100124
rect 35836 100064 35900 100068
rect 66316 100124 66380 100128
rect 66316 100068 66320 100124
rect 66320 100068 66376 100124
rect 66376 100068 66380 100124
rect 66316 100064 66380 100068
rect 66396 100124 66460 100128
rect 66396 100068 66400 100124
rect 66400 100068 66456 100124
rect 66456 100068 66460 100124
rect 66396 100064 66460 100068
rect 66476 100124 66540 100128
rect 66476 100068 66480 100124
rect 66480 100068 66536 100124
rect 66536 100068 66540 100124
rect 66476 100064 66540 100068
rect 66556 100124 66620 100128
rect 66556 100068 66560 100124
rect 66560 100068 66616 100124
rect 66616 100068 66620 100124
rect 66556 100064 66620 100068
rect 97036 100124 97100 100128
rect 97036 100068 97040 100124
rect 97040 100068 97096 100124
rect 97096 100068 97100 100124
rect 97036 100064 97100 100068
rect 97116 100124 97180 100128
rect 97116 100068 97120 100124
rect 97120 100068 97176 100124
rect 97176 100068 97180 100124
rect 97116 100064 97180 100068
rect 97196 100124 97260 100128
rect 97196 100068 97200 100124
rect 97200 100068 97256 100124
rect 97256 100068 97260 100124
rect 97196 100064 97260 100068
rect 97276 100124 97340 100128
rect 97276 100068 97280 100124
rect 97280 100068 97336 100124
rect 97336 100068 97340 100124
rect 97276 100064 97340 100068
rect 4216 99580 4280 99584
rect 4216 99524 4220 99580
rect 4220 99524 4276 99580
rect 4276 99524 4280 99580
rect 4216 99520 4280 99524
rect 4296 99580 4360 99584
rect 4296 99524 4300 99580
rect 4300 99524 4356 99580
rect 4356 99524 4360 99580
rect 4296 99520 4360 99524
rect 4376 99580 4440 99584
rect 4376 99524 4380 99580
rect 4380 99524 4436 99580
rect 4436 99524 4440 99580
rect 4376 99520 4440 99524
rect 4456 99580 4520 99584
rect 4456 99524 4460 99580
rect 4460 99524 4516 99580
rect 4516 99524 4520 99580
rect 4456 99520 4520 99524
rect 34936 99580 35000 99584
rect 34936 99524 34940 99580
rect 34940 99524 34996 99580
rect 34996 99524 35000 99580
rect 34936 99520 35000 99524
rect 35016 99580 35080 99584
rect 35016 99524 35020 99580
rect 35020 99524 35076 99580
rect 35076 99524 35080 99580
rect 35016 99520 35080 99524
rect 35096 99580 35160 99584
rect 35096 99524 35100 99580
rect 35100 99524 35156 99580
rect 35156 99524 35160 99580
rect 35096 99520 35160 99524
rect 35176 99580 35240 99584
rect 35176 99524 35180 99580
rect 35180 99524 35236 99580
rect 35236 99524 35240 99580
rect 35176 99520 35240 99524
rect 65656 99580 65720 99584
rect 65656 99524 65660 99580
rect 65660 99524 65716 99580
rect 65716 99524 65720 99580
rect 65656 99520 65720 99524
rect 65736 99580 65800 99584
rect 65736 99524 65740 99580
rect 65740 99524 65796 99580
rect 65796 99524 65800 99580
rect 65736 99520 65800 99524
rect 65816 99580 65880 99584
rect 65816 99524 65820 99580
rect 65820 99524 65876 99580
rect 65876 99524 65880 99580
rect 65816 99520 65880 99524
rect 65896 99580 65960 99584
rect 65896 99524 65900 99580
rect 65900 99524 65956 99580
rect 65956 99524 65960 99580
rect 65896 99520 65960 99524
rect 96376 99580 96440 99584
rect 96376 99524 96380 99580
rect 96380 99524 96436 99580
rect 96436 99524 96440 99580
rect 96376 99520 96440 99524
rect 96456 99580 96520 99584
rect 96456 99524 96460 99580
rect 96460 99524 96516 99580
rect 96516 99524 96520 99580
rect 96456 99520 96520 99524
rect 96536 99580 96600 99584
rect 96536 99524 96540 99580
rect 96540 99524 96596 99580
rect 96596 99524 96600 99580
rect 96536 99520 96600 99524
rect 96616 99580 96680 99584
rect 96616 99524 96620 99580
rect 96620 99524 96676 99580
rect 96676 99524 96680 99580
rect 96616 99520 96680 99524
rect 4876 99036 4940 99040
rect 4876 98980 4880 99036
rect 4880 98980 4936 99036
rect 4936 98980 4940 99036
rect 4876 98976 4940 98980
rect 4956 99036 5020 99040
rect 4956 98980 4960 99036
rect 4960 98980 5016 99036
rect 5016 98980 5020 99036
rect 4956 98976 5020 98980
rect 5036 99036 5100 99040
rect 5036 98980 5040 99036
rect 5040 98980 5096 99036
rect 5096 98980 5100 99036
rect 5036 98976 5100 98980
rect 5116 99036 5180 99040
rect 5116 98980 5120 99036
rect 5120 98980 5176 99036
rect 5176 98980 5180 99036
rect 5116 98976 5180 98980
rect 35596 99036 35660 99040
rect 35596 98980 35600 99036
rect 35600 98980 35656 99036
rect 35656 98980 35660 99036
rect 35596 98976 35660 98980
rect 35676 99036 35740 99040
rect 35676 98980 35680 99036
rect 35680 98980 35736 99036
rect 35736 98980 35740 99036
rect 35676 98976 35740 98980
rect 35756 99036 35820 99040
rect 35756 98980 35760 99036
rect 35760 98980 35816 99036
rect 35816 98980 35820 99036
rect 35756 98976 35820 98980
rect 35836 99036 35900 99040
rect 35836 98980 35840 99036
rect 35840 98980 35896 99036
rect 35896 98980 35900 99036
rect 35836 98976 35900 98980
rect 66316 99036 66380 99040
rect 66316 98980 66320 99036
rect 66320 98980 66376 99036
rect 66376 98980 66380 99036
rect 66316 98976 66380 98980
rect 66396 99036 66460 99040
rect 66396 98980 66400 99036
rect 66400 98980 66456 99036
rect 66456 98980 66460 99036
rect 66396 98976 66460 98980
rect 66476 99036 66540 99040
rect 66476 98980 66480 99036
rect 66480 98980 66536 99036
rect 66536 98980 66540 99036
rect 66476 98976 66540 98980
rect 66556 99036 66620 99040
rect 66556 98980 66560 99036
rect 66560 98980 66616 99036
rect 66616 98980 66620 99036
rect 66556 98976 66620 98980
rect 97036 99036 97100 99040
rect 97036 98980 97040 99036
rect 97040 98980 97096 99036
rect 97096 98980 97100 99036
rect 97036 98976 97100 98980
rect 97116 99036 97180 99040
rect 97116 98980 97120 99036
rect 97120 98980 97176 99036
rect 97176 98980 97180 99036
rect 97116 98976 97180 98980
rect 97196 99036 97260 99040
rect 97196 98980 97200 99036
rect 97200 98980 97256 99036
rect 97256 98980 97260 99036
rect 97196 98976 97260 98980
rect 97276 99036 97340 99040
rect 97276 98980 97280 99036
rect 97280 98980 97336 99036
rect 97336 98980 97340 99036
rect 97276 98976 97340 98980
rect 4216 98492 4280 98496
rect 4216 98436 4220 98492
rect 4220 98436 4276 98492
rect 4276 98436 4280 98492
rect 4216 98432 4280 98436
rect 4296 98492 4360 98496
rect 4296 98436 4300 98492
rect 4300 98436 4356 98492
rect 4356 98436 4360 98492
rect 4296 98432 4360 98436
rect 4376 98492 4440 98496
rect 4376 98436 4380 98492
rect 4380 98436 4436 98492
rect 4436 98436 4440 98492
rect 4376 98432 4440 98436
rect 4456 98492 4520 98496
rect 4456 98436 4460 98492
rect 4460 98436 4516 98492
rect 4516 98436 4520 98492
rect 4456 98432 4520 98436
rect 34936 98492 35000 98496
rect 34936 98436 34940 98492
rect 34940 98436 34996 98492
rect 34996 98436 35000 98492
rect 34936 98432 35000 98436
rect 35016 98492 35080 98496
rect 35016 98436 35020 98492
rect 35020 98436 35076 98492
rect 35076 98436 35080 98492
rect 35016 98432 35080 98436
rect 35096 98492 35160 98496
rect 35096 98436 35100 98492
rect 35100 98436 35156 98492
rect 35156 98436 35160 98492
rect 35096 98432 35160 98436
rect 35176 98492 35240 98496
rect 35176 98436 35180 98492
rect 35180 98436 35236 98492
rect 35236 98436 35240 98492
rect 35176 98432 35240 98436
rect 65656 98492 65720 98496
rect 65656 98436 65660 98492
rect 65660 98436 65716 98492
rect 65716 98436 65720 98492
rect 65656 98432 65720 98436
rect 65736 98492 65800 98496
rect 65736 98436 65740 98492
rect 65740 98436 65796 98492
rect 65796 98436 65800 98492
rect 65736 98432 65800 98436
rect 65816 98492 65880 98496
rect 65816 98436 65820 98492
rect 65820 98436 65876 98492
rect 65876 98436 65880 98492
rect 65816 98432 65880 98436
rect 65896 98492 65960 98496
rect 65896 98436 65900 98492
rect 65900 98436 65956 98492
rect 65956 98436 65960 98492
rect 65896 98432 65960 98436
rect 96376 98492 96440 98496
rect 96376 98436 96380 98492
rect 96380 98436 96436 98492
rect 96436 98436 96440 98492
rect 96376 98432 96440 98436
rect 96456 98492 96520 98496
rect 96456 98436 96460 98492
rect 96460 98436 96516 98492
rect 96516 98436 96520 98492
rect 96456 98432 96520 98436
rect 96536 98492 96600 98496
rect 96536 98436 96540 98492
rect 96540 98436 96596 98492
rect 96596 98436 96600 98492
rect 96536 98432 96600 98436
rect 96616 98492 96680 98496
rect 96616 98436 96620 98492
rect 96620 98436 96676 98492
rect 96676 98436 96680 98492
rect 96616 98432 96680 98436
rect 4876 97948 4940 97952
rect 4876 97892 4880 97948
rect 4880 97892 4936 97948
rect 4936 97892 4940 97948
rect 4876 97888 4940 97892
rect 4956 97948 5020 97952
rect 4956 97892 4960 97948
rect 4960 97892 5016 97948
rect 5016 97892 5020 97948
rect 4956 97888 5020 97892
rect 5036 97948 5100 97952
rect 5036 97892 5040 97948
rect 5040 97892 5096 97948
rect 5096 97892 5100 97948
rect 5036 97888 5100 97892
rect 5116 97948 5180 97952
rect 5116 97892 5120 97948
rect 5120 97892 5176 97948
rect 5176 97892 5180 97948
rect 5116 97888 5180 97892
rect 35596 97948 35660 97952
rect 35596 97892 35600 97948
rect 35600 97892 35656 97948
rect 35656 97892 35660 97948
rect 35596 97888 35660 97892
rect 35676 97948 35740 97952
rect 35676 97892 35680 97948
rect 35680 97892 35736 97948
rect 35736 97892 35740 97948
rect 35676 97888 35740 97892
rect 35756 97948 35820 97952
rect 35756 97892 35760 97948
rect 35760 97892 35816 97948
rect 35816 97892 35820 97948
rect 35756 97888 35820 97892
rect 35836 97948 35900 97952
rect 35836 97892 35840 97948
rect 35840 97892 35896 97948
rect 35896 97892 35900 97948
rect 35836 97888 35900 97892
rect 66316 97948 66380 97952
rect 66316 97892 66320 97948
rect 66320 97892 66376 97948
rect 66376 97892 66380 97948
rect 66316 97888 66380 97892
rect 66396 97948 66460 97952
rect 66396 97892 66400 97948
rect 66400 97892 66456 97948
rect 66456 97892 66460 97948
rect 66396 97888 66460 97892
rect 66476 97948 66540 97952
rect 66476 97892 66480 97948
rect 66480 97892 66536 97948
rect 66536 97892 66540 97948
rect 66476 97888 66540 97892
rect 66556 97948 66620 97952
rect 66556 97892 66560 97948
rect 66560 97892 66616 97948
rect 66616 97892 66620 97948
rect 66556 97888 66620 97892
rect 97036 97948 97100 97952
rect 97036 97892 97040 97948
rect 97040 97892 97096 97948
rect 97096 97892 97100 97948
rect 97036 97888 97100 97892
rect 97116 97948 97180 97952
rect 97116 97892 97120 97948
rect 97120 97892 97176 97948
rect 97176 97892 97180 97948
rect 97116 97888 97180 97892
rect 97196 97948 97260 97952
rect 97196 97892 97200 97948
rect 97200 97892 97256 97948
rect 97256 97892 97260 97948
rect 97196 97888 97260 97892
rect 97276 97948 97340 97952
rect 97276 97892 97280 97948
rect 97280 97892 97336 97948
rect 97336 97892 97340 97948
rect 97276 97888 97340 97892
rect 4216 97404 4280 97408
rect 4216 97348 4220 97404
rect 4220 97348 4276 97404
rect 4276 97348 4280 97404
rect 4216 97344 4280 97348
rect 4296 97404 4360 97408
rect 4296 97348 4300 97404
rect 4300 97348 4356 97404
rect 4356 97348 4360 97404
rect 4296 97344 4360 97348
rect 4376 97404 4440 97408
rect 4376 97348 4380 97404
rect 4380 97348 4436 97404
rect 4436 97348 4440 97404
rect 4376 97344 4440 97348
rect 4456 97404 4520 97408
rect 4456 97348 4460 97404
rect 4460 97348 4516 97404
rect 4516 97348 4520 97404
rect 4456 97344 4520 97348
rect 34936 97404 35000 97408
rect 34936 97348 34940 97404
rect 34940 97348 34996 97404
rect 34996 97348 35000 97404
rect 34936 97344 35000 97348
rect 35016 97404 35080 97408
rect 35016 97348 35020 97404
rect 35020 97348 35076 97404
rect 35076 97348 35080 97404
rect 35016 97344 35080 97348
rect 35096 97404 35160 97408
rect 35096 97348 35100 97404
rect 35100 97348 35156 97404
rect 35156 97348 35160 97404
rect 35096 97344 35160 97348
rect 35176 97404 35240 97408
rect 35176 97348 35180 97404
rect 35180 97348 35236 97404
rect 35236 97348 35240 97404
rect 35176 97344 35240 97348
rect 65656 97404 65720 97408
rect 65656 97348 65660 97404
rect 65660 97348 65716 97404
rect 65716 97348 65720 97404
rect 65656 97344 65720 97348
rect 65736 97404 65800 97408
rect 65736 97348 65740 97404
rect 65740 97348 65796 97404
rect 65796 97348 65800 97404
rect 65736 97344 65800 97348
rect 65816 97404 65880 97408
rect 65816 97348 65820 97404
rect 65820 97348 65876 97404
rect 65876 97348 65880 97404
rect 65816 97344 65880 97348
rect 65896 97404 65960 97408
rect 65896 97348 65900 97404
rect 65900 97348 65956 97404
rect 65956 97348 65960 97404
rect 65896 97344 65960 97348
rect 96376 97404 96440 97408
rect 96376 97348 96380 97404
rect 96380 97348 96436 97404
rect 96436 97348 96440 97404
rect 96376 97344 96440 97348
rect 96456 97404 96520 97408
rect 96456 97348 96460 97404
rect 96460 97348 96516 97404
rect 96516 97348 96520 97404
rect 96456 97344 96520 97348
rect 96536 97404 96600 97408
rect 96536 97348 96540 97404
rect 96540 97348 96596 97404
rect 96596 97348 96600 97404
rect 96536 97344 96600 97348
rect 96616 97404 96680 97408
rect 96616 97348 96620 97404
rect 96620 97348 96676 97404
rect 96676 97348 96680 97404
rect 96616 97344 96680 97348
rect 4876 96860 4940 96864
rect 4876 96804 4880 96860
rect 4880 96804 4936 96860
rect 4936 96804 4940 96860
rect 4876 96800 4940 96804
rect 4956 96860 5020 96864
rect 4956 96804 4960 96860
rect 4960 96804 5016 96860
rect 5016 96804 5020 96860
rect 4956 96800 5020 96804
rect 5036 96860 5100 96864
rect 5036 96804 5040 96860
rect 5040 96804 5096 96860
rect 5096 96804 5100 96860
rect 5036 96800 5100 96804
rect 5116 96860 5180 96864
rect 5116 96804 5120 96860
rect 5120 96804 5176 96860
rect 5176 96804 5180 96860
rect 5116 96800 5180 96804
rect 35596 96860 35660 96864
rect 35596 96804 35600 96860
rect 35600 96804 35656 96860
rect 35656 96804 35660 96860
rect 35596 96800 35660 96804
rect 35676 96860 35740 96864
rect 35676 96804 35680 96860
rect 35680 96804 35736 96860
rect 35736 96804 35740 96860
rect 35676 96800 35740 96804
rect 35756 96860 35820 96864
rect 35756 96804 35760 96860
rect 35760 96804 35816 96860
rect 35816 96804 35820 96860
rect 35756 96800 35820 96804
rect 35836 96860 35900 96864
rect 35836 96804 35840 96860
rect 35840 96804 35896 96860
rect 35896 96804 35900 96860
rect 35836 96800 35900 96804
rect 66316 96860 66380 96864
rect 66316 96804 66320 96860
rect 66320 96804 66376 96860
rect 66376 96804 66380 96860
rect 66316 96800 66380 96804
rect 66396 96860 66460 96864
rect 66396 96804 66400 96860
rect 66400 96804 66456 96860
rect 66456 96804 66460 96860
rect 66396 96800 66460 96804
rect 66476 96860 66540 96864
rect 66476 96804 66480 96860
rect 66480 96804 66536 96860
rect 66536 96804 66540 96860
rect 66476 96800 66540 96804
rect 66556 96860 66620 96864
rect 66556 96804 66560 96860
rect 66560 96804 66616 96860
rect 66616 96804 66620 96860
rect 66556 96800 66620 96804
rect 97036 96860 97100 96864
rect 97036 96804 97040 96860
rect 97040 96804 97096 96860
rect 97096 96804 97100 96860
rect 97036 96800 97100 96804
rect 97116 96860 97180 96864
rect 97116 96804 97120 96860
rect 97120 96804 97176 96860
rect 97176 96804 97180 96860
rect 97116 96800 97180 96804
rect 97196 96860 97260 96864
rect 97196 96804 97200 96860
rect 97200 96804 97256 96860
rect 97256 96804 97260 96860
rect 97196 96800 97260 96804
rect 97276 96860 97340 96864
rect 97276 96804 97280 96860
rect 97280 96804 97336 96860
rect 97336 96804 97340 96860
rect 97276 96800 97340 96804
rect 4216 96316 4280 96320
rect 4216 96260 4220 96316
rect 4220 96260 4276 96316
rect 4276 96260 4280 96316
rect 4216 96256 4280 96260
rect 4296 96316 4360 96320
rect 4296 96260 4300 96316
rect 4300 96260 4356 96316
rect 4356 96260 4360 96316
rect 4296 96256 4360 96260
rect 4376 96316 4440 96320
rect 4376 96260 4380 96316
rect 4380 96260 4436 96316
rect 4436 96260 4440 96316
rect 4376 96256 4440 96260
rect 4456 96316 4520 96320
rect 4456 96260 4460 96316
rect 4460 96260 4516 96316
rect 4516 96260 4520 96316
rect 4456 96256 4520 96260
rect 34936 96316 35000 96320
rect 34936 96260 34940 96316
rect 34940 96260 34996 96316
rect 34996 96260 35000 96316
rect 34936 96256 35000 96260
rect 35016 96316 35080 96320
rect 35016 96260 35020 96316
rect 35020 96260 35076 96316
rect 35076 96260 35080 96316
rect 35016 96256 35080 96260
rect 35096 96316 35160 96320
rect 35096 96260 35100 96316
rect 35100 96260 35156 96316
rect 35156 96260 35160 96316
rect 35096 96256 35160 96260
rect 35176 96316 35240 96320
rect 35176 96260 35180 96316
rect 35180 96260 35236 96316
rect 35236 96260 35240 96316
rect 35176 96256 35240 96260
rect 65656 96316 65720 96320
rect 65656 96260 65660 96316
rect 65660 96260 65716 96316
rect 65716 96260 65720 96316
rect 65656 96256 65720 96260
rect 65736 96316 65800 96320
rect 65736 96260 65740 96316
rect 65740 96260 65796 96316
rect 65796 96260 65800 96316
rect 65736 96256 65800 96260
rect 65816 96316 65880 96320
rect 65816 96260 65820 96316
rect 65820 96260 65876 96316
rect 65876 96260 65880 96316
rect 65816 96256 65880 96260
rect 65896 96316 65960 96320
rect 65896 96260 65900 96316
rect 65900 96260 65956 96316
rect 65956 96260 65960 96316
rect 65896 96256 65960 96260
rect 96376 96316 96440 96320
rect 96376 96260 96380 96316
rect 96380 96260 96436 96316
rect 96436 96260 96440 96316
rect 96376 96256 96440 96260
rect 96456 96316 96520 96320
rect 96456 96260 96460 96316
rect 96460 96260 96516 96316
rect 96516 96260 96520 96316
rect 96456 96256 96520 96260
rect 96536 96316 96600 96320
rect 96536 96260 96540 96316
rect 96540 96260 96596 96316
rect 96596 96260 96600 96316
rect 96536 96256 96600 96260
rect 96616 96316 96680 96320
rect 96616 96260 96620 96316
rect 96620 96260 96676 96316
rect 96676 96260 96680 96316
rect 96616 96256 96680 96260
rect 4876 95772 4940 95776
rect 4876 95716 4880 95772
rect 4880 95716 4936 95772
rect 4936 95716 4940 95772
rect 4876 95712 4940 95716
rect 4956 95772 5020 95776
rect 4956 95716 4960 95772
rect 4960 95716 5016 95772
rect 5016 95716 5020 95772
rect 4956 95712 5020 95716
rect 5036 95772 5100 95776
rect 5036 95716 5040 95772
rect 5040 95716 5096 95772
rect 5096 95716 5100 95772
rect 5036 95712 5100 95716
rect 5116 95772 5180 95776
rect 5116 95716 5120 95772
rect 5120 95716 5176 95772
rect 5176 95716 5180 95772
rect 5116 95712 5180 95716
rect 35596 95772 35660 95776
rect 35596 95716 35600 95772
rect 35600 95716 35656 95772
rect 35656 95716 35660 95772
rect 35596 95712 35660 95716
rect 35676 95772 35740 95776
rect 35676 95716 35680 95772
rect 35680 95716 35736 95772
rect 35736 95716 35740 95772
rect 35676 95712 35740 95716
rect 35756 95772 35820 95776
rect 35756 95716 35760 95772
rect 35760 95716 35816 95772
rect 35816 95716 35820 95772
rect 35756 95712 35820 95716
rect 35836 95772 35900 95776
rect 35836 95716 35840 95772
rect 35840 95716 35896 95772
rect 35896 95716 35900 95772
rect 35836 95712 35900 95716
rect 66316 95772 66380 95776
rect 66316 95716 66320 95772
rect 66320 95716 66376 95772
rect 66376 95716 66380 95772
rect 66316 95712 66380 95716
rect 66396 95772 66460 95776
rect 66396 95716 66400 95772
rect 66400 95716 66456 95772
rect 66456 95716 66460 95772
rect 66396 95712 66460 95716
rect 66476 95772 66540 95776
rect 66476 95716 66480 95772
rect 66480 95716 66536 95772
rect 66536 95716 66540 95772
rect 66476 95712 66540 95716
rect 66556 95772 66620 95776
rect 66556 95716 66560 95772
rect 66560 95716 66616 95772
rect 66616 95716 66620 95772
rect 66556 95712 66620 95716
rect 97036 95772 97100 95776
rect 97036 95716 97040 95772
rect 97040 95716 97096 95772
rect 97096 95716 97100 95772
rect 97036 95712 97100 95716
rect 97116 95772 97180 95776
rect 97116 95716 97120 95772
rect 97120 95716 97176 95772
rect 97176 95716 97180 95772
rect 97116 95712 97180 95716
rect 97196 95772 97260 95776
rect 97196 95716 97200 95772
rect 97200 95716 97256 95772
rect 97256 95716 97260 95772
rect 97196 95712 97260 95716
rect 97276 95772 97340 95776
rect 97276 95716 97280 95772
rect 97280 95716 97336 95772
rect 97336 95716 97340 95772
rect 97276 95712 97340 95716
rect 4216 95228 4280 95232
rect 4216 95172 4220 95228
rect 4220 95172 4276 95228
rect 4276 95172 4280 95228
rect 4216 95168 4280 95172
rect 4296 95228 4360 95232
rect 4296 95172 4300 95228
rect 4300 95172 4356 95228
rect 4356 95172 4360 95228
rect 4296 95168 4360 95172
rect 4376 95228 4440 95232
rect 4376 95172 4380 95228
rect 4380 95172 4436 95228
rect 4436 95172 4440 95228
rect 4376 95168 4440 95172
rect 4456 95228 4520 95232
rect 4456 95172 4460 95228
rect 4460 95172 4516 95228
rect 4516 95172 4520 95228
rect 4456 95168 4520 95172
rect 34936 95228 35000 95232
rect 34936 95172 34940 95228
rect 34940 95172 34996 95228
rect 34996 95172 35000 95228
rect 34936 95168 35000 95172
rect 35016 95228 35080 95232
rect 35016 95172 35020 95228
rect 35020 95172 35076 95228
rect 35076 95172 35080 95228
rect 35016 95168 35080 95172
rect 35096 95228 35160 95232
rect 35096 95172 35100 95228
rect 35100 95172 35156 95228
rect 35156 95172 35160 95228
rect 35096 95168 35160 95172
rect 35176 95228 35240 95232
rect 35176 95172 35180 95228
rect 35180 95172 35236 95228
rect 35236 95172 35240 95228
rect 35176 95168 35240 95172
rect 65656 95228 65720 95232
rect 65656 95172 65660 95228
rect 65660 95172 65716 95228
rect 65716 95172 65720 95228
rect 65656 95168 65720 95172
rect 65736 95228 65800 95232
rect 65736 95172 65740 95228
rect 65740 95172 65796 95228
rect 65796 95172 65800 95228
rect 65736 95168 65800 95172
rect 65816 95228 65880 95232
rect 65816 95172 65820 95228
rect 65820 95172 65876 95228
rect 65876 95172 65880 95228
rect 65816 95168 65880 95172
rect 65896 95228 65960 95232
rect 65896 95172 65900 95228
rect 65900 95172 65956 95228
rect 65956 95172 65960 95228
rect 65896 95168 65960 95172
rect 96376 95228 96440 95232
rect 96376 95172 96380 95228
rect 96380 95172 96436 95228
rect 96436 95172 96440 95228
rect 96376 95168 96440 95172
rect 96456 95228 96520 95232
rect 96456 95172 96460 95228
rect 96460 95172 96516 95228
rect 96516 95172 96520 95228
rect 96456 95168 96520 95172
rect 96536 95228 96600 95232
rect 96536 95172 96540 95228
rect 96540 95172 96596 95228
rect 96596 95172 96600 95228
rect 96536 95168 96600 95172
rect 96616 95228 96680 95232
rect 96616 95172 96620 95228
rect 96620 95172 96676 95228
rect 96676 95172 96680 95228
rect 96616 95168 96680 95172
rect 4876 94684 4940 94688
rect 4876 94628 4880 94684
rect 4880 94628 4936 94684
rect 4936 94628 4940 94684
rect 4876 94624 4940 94628
rect 4956 94684 5020 94688
rect 4956 94628 4960 94684
rect 4960 94628 5016 94684
rect 5016 94628 5020 94684
rect 4956 94624 5020 94628
rect 5036 94684 5100 94688
rect 5036 94628 5040 94684
rect 5040 94628 5096 94684
rect 5096 94628 5100 94684
rect 5036 94624 5100 94628
rect 5116 94684 5180 94688
rect 5116 94628 5120 94684
rect 5120 94628 5176 94684
rect 5176 94628 5180 94684
rect 5116 94624 5180 94628
rect 35596 94684 35660 94688
rect 35596 94628 35600 94684
rect 35600 94628 35656 94684
rect 35656 94628 35660 94684
rect 35596 94624 35660 94628
rect 35676 94684 35740 94688
rect 35676 94628 35680 94684
rect 35680 94628 35736 94684
rect 35736 94628 35740 94684
rect 35676 94624 35740 94628
rect 35756 94684 35820 94688
rect 35756 94628 35760 94684
rect 35760 94628 35816 94684
rect 35816 94628 35820 94684
rect 35756 94624 35820 94628
rect 35836 94684 35900 94688
rect 35836 94628 35840 94684
rect 35840 94628 35896 94684
rect 35896 94628 35900 94684
rect 35836 94624 35900 94628
rect 66316 94684 66380 94688
rect 66316 94628 66320 94684
rect 66320 94628 66376 94684
rect 66376 94628 66380 94684
rect 66316 94624 66380 94628
rect 66396 94684 66460 94688
rect 66396 94628 66400 94684
rect 66400 94628 66456 94684
rect 66456 94628 66460 94684
rect 66396 94624 66460 94628
rect 66476 94684 66540 94688
rect 66476 94628 66480 94684
rect 66480 94628 66536 94684
rect 66536 94628 66540 94684
rect 66476 94624 66540 94628
rect 66556 94684 66620 94688
rect 66556 94628 66560 94684
rect 66560 94628 66616 94684
rect 66616 94628 66620 94684
rect 66556 94624 66620 94628
rect 97036 94684 97100 94688
rect 97036 94628 97040 94684
rect 97040 94628 97096 94684
rect 97096 94628 97100 94684
rect 97036 94624 97100 94628
rect 97116 94684 97180 94688
rect 97116 94628 97120 94684
rect 97120 94628 97176 94684
rect 97176 94628 97180 94684
rect 97116 94624 97180 94628
rect 97196 94684 97260 94688
rect 97196 94628 97200 94684
rect 97200 94628 97256 94684
rect 97256 94628 97260 94684
rect 97196 94624 97260 94628
rect 97276 94684 97340 94688
rect 97276 94628 97280 94684
rect 97280 94628 97336 94684
rect 97336 94628 97340 94684
rect 97276 94624 97340 94628
rect 4216 94140 4280 94144
rect 4216 94084 4220 94140
rect 4220 94084 4276 94140
rect 4276 94084 4280 94140
rect 4216 94080 4280 94084
rect 4296 94140 4360 94144
rect 4296 94084 4300 94140
rect 4300 94084 4356 94140
rect 4356 94084 4360 94140
rect 4296 94080 4360 94084
rect 4376 94140 4440 94144
rect 4376 94084 4380 94140
rect 4380 94084 4436 94140
rect 4436 94084 4440 94140
rect 4376 94080 4440 94084
rect 4456 94140 4520 94144
rect 4456 94084 4460 94140
rect 4460 94084 4516 94140
rect 4516 94084 4520 94140
rect 4456 94080 4520 94084
rect 34936 94140 35000 94144
rect 34936 94084 34940 94140
rect 34940 94084 34996 94140
rect 34996 94084 35000 94140
rect 34936 94080 35000 94084
rect 35016 94140 35080 94144
rect 35016 94084 35020 94140
rect 35020 94084 35076 94140
rect 35076 94084 35080 94140
rect 35016 94080 35080 94084
rect 35096 94140 35160 94144
rect 35096 94084 35100 94140
rect 35100 94084 35156 94140
rect 35156 94084 35160 94140
rect 35096 94080 35160 94084
rect 35176 94140 35240 94144
rect 35176 94084 35180 94140
rect 35180 94084 35236 94140
rect 35236 94084 35240 94140
rect 35176 94080 35240 94084
rect 65656 94140 65720 94144
rect 65656 94084 65660 94140
rect 65660 94084 65716 94140
rect 65716 94084 65720 94140
rect 65656 94080 65720 94084
rect 65736 94140 65800 94144
rect 65736 94084 65740 94140
rect 65740 94084 65796 94140
rect 65796 94084 65800 94140
rect 65736 94080 65800 94084
rect 65816 94140 65880 94144
rect 65816 94084 65820 94140
rect 65820 94084 65876 94140
rect 65876 94084 65880 94140
rect 65816 94080 65880 94084
rect 65896 94140 65960 94144
rect 65896 94084 65900 94140
rect 65900 94084 65956 94140
rect 65956 94084 65960 94140
rect 65896 94080 65960 94084
rect 96376 94140 96440 94144
rect 96376 94084 96380 94140
rect 96380 94084 96436 94140
rect 96436 94084 96440 94140
rect 96376 94080 96440 94084
rect 96456 94140 96520 94144
rect 96456 94084 96460 94140
rect 96460 94084 96516 94140
rect 96516 94084 96520 94140
rect 96456 94080 96520 94084
rect 96536 94140 96600 94144
rect 96536 94084 96540 94140
rect 96540 94084 96596 94140
rect 96596 94084 96600 94140
rect 96536 94080 96600 94084
rect 96616 94140 96680 94144
rect 96616 94084 96620 94140
rect 96620 94084 96676 94140
rect 96676 94084 96680 94140
rect 96616 94080 96680 94084
rect 4876 93596 4940 93600
rect 4876 93540 4880 93596
rect 4880 93540 4936 93596
rect 4936 93540 4940 93596
rect 4876 93536 4940 93540
rect 4956 93596 5020 93600
rect 4956 93540 4960 93596
rect 4960 93540 5016 93596
rect 5016 93540 5020 93596
rect 4956 93536 5020 93540
rect 5036 93596 5100 93600
rect 5036 93540 5040 93596
rect 5040 93540 5096 93596
rect 5096 93540 5100 93596
rect 5036 93536 5100 93540
rect 5116 93596 5180 93600
rect 5116 93540 5120 93596
rect 5120 93540 5176 93596
rect 5176 93540 5180 93596
rect 5116 93536 5180 93540
rect 35596 93596 35660 93600
rect 35596 93540 35600 93596
rect 35600 93540 35656 93596
rect 35656 93540 35660 93596
rect 35596 93536 35660 93540
rect 35676 93596 35740 93600
rect 35676 93540 35680 93596
rect 35680 93540 35736 93596
rect 35736 93540 35740 93596
rect 35676 93536 35740 93540
rect 35756 93596 35820 93600
rect 35756 93540 35760 93596
rect 35760 93540 35816 93596
rect 35816 93540 35820 93596
rect 35756 93536 35820 93540
rect 35836 93596 35900 93600
rect 35836 93540 35840 93596
rect 35840 93540 35896 93596
rect 35896 93540 35900 93596
rect 35836 93536 35900 93540
rect 66316 93596 66380 93600
rect 66316 93540 66320 93596
rect 66320 93540 66376 93596
rect 66376 93540 66380 93596
rect 66316 93536 66380 93540
rect 66396 93596 66460 93600
rect 66396 93540 66400 93596
rect 66400 93540 66456 93596
rect 66456 93540 66460 93596
rect 66396 93536 66460 93540
rect 66476 93596 66540 93600
rect 66476 93540 66480 93596
rect 66480 93540 66536 93596
rect 66536 93540 66540 93596
rect 66476 93536 66540 93540
rect 66556 93596 66620 93600
rect 66556 93540 66560 93596
rect 66560 93540 66616 93596
rect 66616 93540 66620 93596
rect 66556 93536 66620 93540
rect 97036 93596 97100 93600
rect 97036 93540 97040 93596
rect 97040 93540 97096 93596
rect 97096 93540 97100 93596
rect 97036 93536 97100 93540
rect 97116 93596 97180 93600
rect 97116 93540 97120 93596
rect 97120 93540 97176 93596
rect 97176 93540 97180 93596
rect 97116 93536 97180 93540
rect 97196 93596 97260 93600
rect 97196 93540 97200 93596
rect 97200 93540 97256 93596
rect 97256 93540 97260 93596
rect 97196 93536 97260 93540
rect 97276 93596 97340 93600
rect 97276 93540 97280 93596
rect 97280 93540 97336 93596
rect 97336 93540 97340 93596
rect 97276 93536 97340 93540
rect 4216 93052 4280 93056
rect 4216 92996 4220 93052
rect 4220 92996 4276 93052
rect 4276 92996 4280 93052
rect 4216 92992 4280 92996
rect 4296 93052 4360 93056
rect 4296 92996 4300 93052
rect 4300 92996 4356 93052
rect 4356 92996 4360 93052
rect 4296 92992 4360 92996
rect 4376 93052 4440 93056
rect 4376 92996 4380 93052
rect 4380 92996 4436 93052
rect 4436 92996 4440 93052
rect 4376 92992 4440 92996
rect 4456 93052 4520 93056
rect 4456 92996 4460 93052
rect 4460 92996 4516 93052
rect 4516 92996 4520 93052
rect 4456 92992 4520 92996
rect 34936 93052 35000 93056
rect 34936 92996 34940 93052
rect 34940 92996 34996 93052
rect 34996 92996 35000 93052
rect 34936 92992 35000 92996
rect 35016 93052 35080 93056
rect 35016 92996 35020 93052
rect 35020 92996 35076 93052
rect 35076 92996 35080 93052
rect 35016 92992 35080 92996
rect 35096 93052 35160 93056
rect 35096 92996 35100 93052
rect 35100 92996 35156 93052
rect 35156 92996 35160 93052
rect 35096 92992 35160 92996
rect 35176 93052 35240 93056
rect 35176 92996 35180 93052
rect 35180 92996 35236 93052
rect 35236 92996 35240 93052
rect 35176 92992 35240 92996
rect 65656 93052 65720 93056
rect 65656 92996 65660 93052
rect 65660 92996 65716 93052
rect 65716 92996 65720 93052
rect 65656 92992 65720 92996
rect 65736 93052 65800 93056
rect 65736 92996 65740 93052
rect 65740 92996 65796 93052
rect 65796 92996 65800 93052
rect 65736 92992 65800 92996
rect 65816 93052 65880 93056
rect 65816 92996 65820 93052
rect 65820 92996 65876 93052
rect 65876 92996 65880 93052
rect 65816 92992 65880 92996
rect 65896 93052 65960 93056
rect 65896 92996 65900 93052
rect 65900 92996 65956 93052
rect 65956 92996 65960 93052
rect 65896 92992 65960 92996
rect 96376 93052 96440 93056
rect 96376 92996 96380 93052
rect 96380 92996 96436 93052
rect 96436 92996 96440 93052
rect 96376 92992 96440 92996
rect 96456 93052 96520 93056
rect 96456 92996 96460 93052
rect 96460 92996 96516 93052
rect 96516 92996 96520 93052
rect 96456 92992 96520 92996
rect 96536 93052 96600 93056
rect 96536 92996 96540 93052
rect 96540 92996 96596 93052
rect 96596 92996 96600 93052
rect 96536 92992 96600 92996
rect 96616 93052 96680 93056
rect 96616 92996 96620 93052
rect 96620 92996 96676 93052
rect 96676 92996 96680 93052
rect 96616 92992 96680 92996
rect 4876 92508 4940 92512
rect 4876 92452 4880 92508
rect 4880 92452 4936 92508
rect 4936 92452 4940 92508
rect 4876 92448 4940 92452
rect 4956 92508 5020 92512
rect 4956 92452 4960 92508
rect 4960 92452 5016 92508
rect 5016 92452 5020 92508
rect 4956 92448 5020 92452
rect 5036 92508 5100 92512
rect 5036 92452 5040 92508
rect 5040 92452 5096 92508
rect 5096 92452 5100 92508
rect 5036 92448 5100 92452
rect 5116 92508 5180 92512
rect 5116 92452 5120 92508
rect 5120 92452 5176 92508
rect 5176 92452 5180 92508
rect 5116 92448 5180 92452
rect 35596 92508 35660 92512
rect 35596 92452 35600 92508
rect 35600 92452 35656 92508
rect 35656 92452 35660 92508
rect 35596 92448 35660 92452
rect 35676 92508 35740 92512
rect 35676 92452 35680 92508
rect 35680 92452 35736 92508
rect 35736 92452 35740 92508
rect 35676 92448 35740 92452
rect 35756 92508 35820 92512
rect 35756 92452 35760 92508
rect 35760 92452 35816 92508
rect 35816 92452 35820 92508
rect 35756 92448 35820 92452
rect 35836 92508 35900 92512
rect 35836 92452 35840 92508
rect 35840 92452 35896 92508
rect 35896 92452 35900 92508
rect 35836 92448 35900 92452
rect 66316 92508 66380 92512
rect 66316 92452 66320 92508
rect 66320 92452 66376 92508
rect 66376 92452 66380 92508
rect 66316 92448 66380 92452
rect 66396 92508 66460 92512
rect 66396 92452 66400 92508
rect 66400 92452 66456 92508
rect 66456 92452 66460 92508
rect 66396 92448 66460 92452
rect 66476 92508 66540 92512
rect 66476 92452 66480 92508
rect 66480 92452 66536 92508
rect 66536 92452 66540 92508
rect 66476 92448 66540 92452
rect 66556 92508 66620 92512
rect 66556 92452 66560 92508
rect 66560 92452 66616 92508
rect 66616 92452 66620 92508
rect 66556 92448 66620 92452
rect 97036 92508 97100 92512
rect 97036 92452 97040 92508
rect 97040 92452 97096 92508
rect 97096 92452 97100 92508
rect 97036 92448 97100 92452
rect 97116 92508 97180 92512
rect 97116 92452 97120 92508
rect 97120 92452 97176 92508
rect 97176 92452 97180 92508
rect 97116 92448 97180 92452
rect 97196 92508 97260 92512
rect 97196 92452 97200 92508
rect 97200 92452 97256 92508
rect 97256 92452 97260 92508
rect 97196 92448 97260 92452
rect 97276 92508 97340 92512
rect 97276 92452 97280 92508
rect 97280 92452 97336 92508
rect 97336 92452 97340 92508
rect 97276 92448 97340 92452
rect 4216 91964 4280 91968
rect 4216 91908 4220 91964
rect 4220 91908 4276 91964
rect 4276 91908 4280 91964
rect 4216 91904 4280 91908
rect 4296 91964 4360 91968
rect 4296 91908 4300 91964
rect 4300 91908 4356 91964
rect 4356 91908 4360 91964
rect 4296 91904 4360 91908
rect 4376 91964 4440 91968
rect 4376 91908 4380 91964
rect 4380 91908 4436 91964
rect 4436 91908 4440 91964
rect 4376 91904 4440 91908
rect 4456 91964 4520 91968
rect 4456 91908 4460 91964
rect 4460 91908 4516 91964
rect 4516 91908 4520 91964
rect 4456 91904 4520 91908
rect 34936 91964 35000 91968
rect 34936 91908 34940 91964
rect 34940 91908 34996 91964
rect 34996 91908 35000 91964
rect 34936 91904 35000 91908
rect 35016 91964 35080 91968
rect 35016 91908 35020 91964
rect 35020 91908 35076 91964
rect 35076 91908 35080 91964
rect 35016 91904 35080 91908
rect 35096 91964 35160 91968
rect 35096 91908 35100 91964
rect 35100 91908 35156 91964
rect 35156 91908 35160 91964
rect 35096 91904 35160 91908
rect 35176 91964 35240 91968
rect 35176 91908 35180 91964
rect 35180 91908 35236 91964
rect 35236 91908 35240 91964
rect 35176 91904 35240 91908
rect 65656 91964 65720 91968
rect 65656 91908 65660 91964
rect 65660 91908 65716 91964
rect 65716 91908 65720 91964
rect 65656 91904 65720 91908
rect 65736 91964 65800 91968
rect 65736 91908 65740 91964
rect 65740 91908 65796 91964
rect 65796 91908 65800 91964
rect 65736 91904 65800 91908
rect 65816 91964 65880 91968
rect 65816 91908 65820 91964
rect 65820 91908 65876 91964
rect 65876 91908 65880 91964
rect 65816 91904 65880 91908
rect 65896 91964 65960 91968
rect 65896 91908 65900 91964
rect 65900 91908 65956 91964
rect 65956 91908 65960 91964
rect 65896 91904 65960 91908
rect 96376 91964 96440 91968
rect 96376 91908 96380 91964
rect 96380 91908 96436 91964
rect 96436 91908 96440 91964
rect 96376 91904 96440 91908
rect 96456 91964 96520 91968
rect 96456 91908 96460 91964
rect 96460 91908 96516 91964
rect 96516 91908 96520 91964
rect 96456 91904 96520 91908
rect 96536 91964 96600 91968
rect 96536 91908 96540 91964
rect 96540 91908 96596 91964
rect 96596 91908 96600 91964
rect 96536 91904 96600 91908
rect 96616 91964 96680 91968
rect 96616 91908 96620 91964
rect 96620 91908 96676 91964
rect 96676 91908 96680 91964
rect 96616 91904 96680 91908
rect 4876 91420 4940 91424
rect 4876 91364 4880 91420
rect 4880 91364 4936 91420
rect 4936 91364 4940 91420
rect 4876 91360 4940 91364
rect 4956 91420 5020 91424
rect 4956 91364 4960 91420
rect 4960 91364 5016 91420
rect 5016 91364 5020 91420
rect 4956 91360 5020 91364
rect 5036 91420 5100 91424
rect 5036 91364 5040 91420
rect 5040 91364 5096 91420
rect 5096 91364 5100 91420
rect 5036 91360 5100 91364
rect 5116 91420 5180 91424
rect 5116 91364 5120 91420
rect 5120 91364 5176 91420
rect 5176 91364 5180 91420
rect 5116 91360 5180 91364
rect 35596 91420 35660 91424
rect 35596 91364 35600 91420
rect 35600 91364 35656 91420
rect 35656 91364 35660 91420
rect 35596 91360 35660 91364
rect 35676 91420 35740 91424
rect 35676 91364 35680 91420
rect 35680 91364 35736 91420
rect 35736 91364 35740 91420
rect 35676 91360 35740 91364
rect 35756 91420 35820 91424
rect 35756 91364 35760 91420
rect 35760 91364 35816 91420
rect 35816 91364 35820 91420
rect 35756 91360 35820 91364
rect 35836 91420 35900 91424
rect 35836 91364 35840 91420
rect 35840 91364 35896 91420
rect 35896 91364 35900 91420
rect 35836 91360 35900 91364
rect 66316 91420 66380 91424
rect 66316 91364 66320 91420
rect 66320 91364 66376 91420
rect 66376 91364 66380 91420
rect 66316 91360 66380 91364
rect 66396 91420 66460 91424
rect 66396 91364 66400 91420
rect 66400 91364 66456 91420
rect 66456 91364 66460 91420
rect 66396 91360 66460 91364
rect 66476 91420 66540 91424
rect 66476 91364 66480 91420
rect 66480 91364 66536 91420
rect 66536 91364 66540 91420
rect 66476 91360 66540 91364
rect 66556 91420 66620 91424
rect 66556 91364 66560 91420
rect 66560 91364 66616 91420
rect 66616 91364 66620 91420
rect 66556 91360 66620 91364
rect 97036 91420 97100 91424
rect 97036 91364 97040 91420
rect 97040 91364 97096 91420
rect 97096 91364 97100 91420
rect 97036 91360 97100 91364
rect 97116 91420 97180 91424
rect 97116 91364 97120 91420
rect 97120 91364 97176 91420
rect 97176 91364 97180 91420
rect 97116 91360 97180 91364
rect 97196 91420 97260 91424
rect 97196 91364 97200 91420
rect 97200 91364 97256 91420
rect 97256 91364 97260 91420
rect 97196 91360 97260 91364
rect 97276 91420 97340 91424
rect 97276 91364 97280 91420
rect 97280 91364 97336 91420
rect 97336 91364 97340 91420
rect 97276 91360 97340 91364
rect 4216 90876 4280 90880
rect 4216 90820 4220 90876
rect 4220 90820 4276 90876
rect 4276 90820 4280 90876
rect 4216 90816 4280 90820
rect 4296 90876 4360 90880
rect 4296 90820 4300 90876
rect 4300 90820 4356 90876
rect 4356 90820 4360 90876
rect 4296 90816 4360 90820
rect 4376 90876 4440 90880
rect 4376 90820 4380 90876
rect 4380 90820 4436 90876
rect 4436 90820 4440 90876
rect 4376 90816 4440 90820
rect 4456 90876 4520 90880
rect 4456 90820 4460 90876
rect 4460 90820 4516 90876
rect 4516 90820 4520 90876
rect 4456 90816 4520 90820
rect 34936 90876 35000 90880
rect 34936 90820 34940 90876
rect 34940 90820 34996 90876
rect 34996 90820 35000 90876
rect 34936 90816 35000 90820
rect 35016 90876 35080 90880
rect 35016 90820 35020 90876
rect 35020 90820 35076 90876
rect 35076 90820 35080 90876
rect 35016 90816 35080 90820
rect 35096 90876 35160 90880
rect 35096 90820 35100 90876
rect 35100 90820 35156 90876
rect 35156 90820 35160 90876
rect 35096 90816 35160 90820
rect 35176 90876 35240 90880
rect 35176 90820 35180 90876
rect 35180 90820 35236 90876
rect 35236 90820 35240 90876
rect 35176 90816 35240 90820
rect 65656 90876 65720 90880
rect 65656 90820 65660 90876
rect 65660 90820 65716 90876
rect 65716 90820 65720 90876
rect 65656 90816 65720 90820
rect 65736 90876 65800 90880
rect 65736 90820 65740 90876
rect 65740 90820 65796 90876
rect 65796 90820 65800 90876
rect 65736 90816 65800 90820
rect 65816 90876 65880 90880
rect 65816 90820 65820 90876
rect 65820 90820 65876 90876
rect 65876 90820 65880 90876
rect 65816 90816 65880 90820
rect 65896 90876 65960 90880
rect 65896 90820 65900 90876
rect 65900 90820 65956 90876
rect 65956 90820 65960 90876
rect 65896 90816 65960 90820
rect 96376 90876 96440 90880
rect 96376 90820 96380 90876
rect 96380 90820 96436 90876
rect 96436 90820 96440 90876
rect 96376 90816 96440 90820
rect 96456 90876 96520 90880
rect 96456 90820 96460 90876
rect 96460 90820 96516 90876
rect 96516 90820 96520 90876
rect 96456 90816 96520 90820
rect 96536 90876 96600 90880
rect 96536 90820 96540 90876
rect 96540 90820 96596 90876
rect 96596 90820 96600 90876
rect 96536 90816 96600 90820
rect 96616 90876 96680 90880
rect 96616 90820 96620 90876
rect 96620 90820 96676 90876
rect 96676 90820 96680 90876
rect 96616 90816 96680 90820
rect 4876 90332 4940 90336
rect 4876 90276 4880 90332
rect 4880 90276 4936 90332
rect 4936 90276 4940 90332
rect 4876 90272 4940 90276
rect 4956 90332 5020 90336
rect 4956 90276 4960 90332
rect 4960 90276 5016 90332
rect 5016 90276 5020 90332
rect 4956 90272 5020 90276
rect 5036 90332 5100 90336
rect 5036 90276 5040 90332
rect 5040 90276 5096 90332
rect 5096 90276 5100 90332
rect 5036 90272 5100 90276
rect 5116 90332 5180 90336
rect 5116 90276 5120 90332
rect 5120 90276 5176 90332
rect 5176 90276 5180 90332
rect 5116 90272 5180 90276
rect 35596 90332 35660 90336
rect 35596 90276 35600 90332
rect 35600 90276 35656 90332
rect 35656 90276 35660 90332
rect 35596 90272 35660 90276
rect 35676 90332 35740 90336
rect 35676 90276 35680 90332
rect 35680 90276 35736 90332
rect 35736 90276 35740 90332
rect 35676 90272 35740 90276
rect 35756 90332 35820 90336
rect 35756 90276 35760 90332
rect 35760 90276 35816 90332
rect 35816 90276 35820 90332
rect 35756 90272 35820 90276
rect 35836 90332 35900 90336
rect 35836 90276 35840 90332
rect 35840 90276 35896 90332
rect 35896 90276 35900 90332
rect 35836 90272 35900 90276
rect 66316 90332 66380 90336
rect 66316 90276 66320 90332
rect 66320 90276 66376 90332
rect 66376 90276 66380 90332
rect 66316 90272 66380 90276
rect 66396 90332 66460 90336
rect 66396 90276 66400 90332
rect 66400 90276 66456 90332
rect 66456 90276 66460 90332
rect 66396 90272 66460 90276
rect 66476 90332 66540 90336
rect 66476 90276 66480 90332
rect 66480 90276 66536 90332
rect 66536 90276 66540 90332
rect 66476 90272 66540 90276
rect 66556 90332 66620 90336
rect 66556 90276 66560 90332
rect 66560 90276 66616 90332
rect 66616 90276 66620 90332
rect 66556 90272 66620 90276
rect 97036 90332 97100 90336
rect 97036 90276 97040 90332
rect 97040 90276 97096 90332
rect 97096 90276 97100 90332
rect 97036 90272 97100 90276
rect 97116 90332 97180 90336
rect 97116 90276 97120 90332
rect 97120 90276 97176 90332
rect 97176 90276 97180 90332
rect 97116 90272 97180 90276
rect 97196 90332 97260 90336
rect 97196 90276 97200 90332
rect 97200 90276 97256 90332
rect 97256 90276 97260 90332
rect 97196 90272 97260 90276
rect 97276 90332 97340 90336
rect 97276 90276 97280 90332
rect 97280 90276 97336 90332
rect 97336 90276 97340 90332
rect 97276 90272 97340 90276
rect 4216 89788 4280 89792
rect 4216 89732 4220 89788
rect 4220 89732 4276 89788
rect 4276 89732 4280 89788
rect 4216 89728 4280 89732
rect 4296 89788 4360 89792
rect 4296 89732 4300 89788
rect 4300 89732 4356 89788
rect 4356 89732 4360 89788
rect 4296 89728 4360 89732
rect 4376 89788 4440 89792
rect 4376 89732 4380 89788
rect 4380 89732 4436 89788
rect 4436 89732 4440 89788
rect 4376 89728 4440 89732
rect 4456 89788 4520 89792
rect 4456 89732 4460 89788
rect 4460 89732 4516 89788
rect 4516 89732 4520 89788
rect 4456 89728 4520 89732
rect 34936 89788 35000 89792
rect 34936 89732 34940 89788
rect 34940 89732 34996 89788
rect 34996 89732 35000 89788
rect 34936 89728 35000 89732
rect 35016 89788 35080 89792
rect 35016 89732 35020 89788
rect 35020 89732 35076 89788
rect 35076 89732 35080 89788
rect 35016 89728 35080 89732
rect 35096 89788 35160 89792
rect 35096 89732 35100 89788
rect 35100 89732 35156 89788
rect 35156 89732 35160 89788
rect 35096 89728 35160 89732
rect 35176 89788 35240 89792
rect 35176 89732 35180 89788
rect 35180 89732 35236 89788
rect 35236 89732 35240 89788
rect 35176 89728 35240 89732
rect 65656 89788 65720 89792
rect 65656 89732 65660 89788
rect 65660 89732 65716 89788
rect 65716 89732 65720 89788
rect 65656 89728 65720 89732
rect 65736 89788 65800 89792
rect 65736 89732 65740 89788
rect 65740 89732 65796 89788
rect 65796 89732 65800 89788
rect 65736 89728 65800 89732
rect 65816 89788 65880 89792
rect 65816 89732 65820 89788
rect 65820 89732 65876 89788
rect 65876 89732 65880 89788
rect 65816 89728 65880 89732
rect 65896 89788 65960 89792
rect 65896 89732 65900 89788
rect 65900 89732 65956 89788
rect 65956 89732 65960 89788
rect 65896 89728 65960 89732
rect 96376 89788 96440 89792
rect 96376 89732 96380 89788
rect 96380 89732 96436 89788
rect 96436 89732 96440 89788
rect 96376 89728 96440 89732
rect 96456 89788 96520 89792
rect 96456 89732 96460 89788
rect 96460 89732 96516 89788
rect 96516 89732 96520 89788
rect 96456 89728 96520 89732
rect 96536 89788 96600 89792
rect 96536 89732 96540 89788
rect 96540 89732 96596 89788
rect 96596 89732 96600 89788
rect 96536 89728 96600 89732
rect 96616 89788 96680 89792
rect 96616 89732 96620 89788
rect 96620 89732 96676 89788
rect 96676 89732 96680 89788
rect 96616 89728 96680 89732
rect 4876 89244 4940 89248
rect 4876 89188 4880 89244
rect 4880 89188 4936 89244
rect 4936 89188 4940 89244
rect 4876 89184 4940 89188
rect 4956 89244 5020 89248
rect 4956 89188 4960 89244
rect 4960 89188 5016 89244
rect 5016 89188 5020 89244
rect 4956 89184 5020 89188
rect 5036 89244 5100 89248
rect 5036 89188 5040 89244
rect 5040 89188 5096 89244
rect 5096 89188 5100 89244
rect 5036 89184 5100 89188
rect 5116 89244 5180 89248
rect 5116 89188 5120 89244
rect 5120 89188 5176 89244
rect 5176 89188 5180 89244
rect 5116 89184 5180 89188
rect 35596 89244 35660 89248
rect 35596 89188 35600 89244
rect 35600 89188 35656 89244
rect 35656 89188 35660 89244
rect 35596 89184 35660 89188
rect 35676 89244 35740 89248
rect 35676 89188 35680 89244
rect 35680 89188 35736 89244
rect 35736 89188 35740 89244
rect 35676 89184 35740 89188
rect 35756 89244 35820 89248
rect 35756 89188 35760 89244
rect 35760 89188 35816 89244
rect 35816 89188 35820 89244
rect 35756 89184 35820 89188
rect 35836 89244 35900 89248
rect 35836 89188 35840 89244
rect 35840 89188 35896 89244
rect 35896 89188 35900 89244
rect 35836 89184 35900 89188
rect 66316 89244 66380 89248
rect 66316 89188 66320 89244
rect 66320 89188 66376 89244
rect 66376 89188 66380 89244
rect 66316 89184 66380 89188
rect 66396 89244 66460 89248
rect 66396 89188 66400 89244
rect 66400 89188 66456 89244
rect 66456 89188 66460 89244
rect 66396 89184 66460 89188
rect 66476 89244 66540 89248
rect 66476 89188 66480 89244
rect 66480 89188 66536 89244
rect 66536 89188 66540 89244
rect 66476 89184 66540 89188
rect 66556 89244 66620 89248
rect 66556 89188 66560 89244
rect 66560 89188 66616 89244
rect 66616 89188 66620 89244
rect 66556 89184 66620 89188
rect 97036 89244 97100 89248
rect 97036 89188 97040 89244
rect 97040 89188 97096 89244
rect 97096 89188 97100 89244
rect 97036 89184 97100 89188
rect 97116 89244 97180 89248
rect 97116 89188 97120 89244
rect 97120 89188 97176 89244
rect 97176 89188 97180 89244
rect 97116 89184 97180 89188
rect 97196 89244 97260 89248
rect 97196 89188 97200 89244
rect 97200 89188 97256 89244
rect 97256 89188 97260 89244
rect 97196 89184 97260 89188
rect 97276 89244 97340 89248
rect 97276 89188 97280 89244
rect 97280 89188 97336 89244
rect 97336 89188 97340 89244
rect 97276 89184 97340 89188
rect 4216 88700 4280 88704
rect 4216 88644 4220 88700
rect 4220 88644 4276 88700
rect 4276 88644 4280 88700
rect 4216 88640 4280 88644
rect 4296 88700 4360 88704
rect 4296 88644 4300 88700
rect 4300 88644 4356 88700
rect 4356 88644 4360 88700
rect 4296 88640 4360 88644
rect 4376 88700 4440 88704
rect 4376 88644 4380 88700
rect 4380 88644 4436 88700
rect 4436 88644 4440 88700
rect 4376 88640 4440 88644
rect 4456 88700 4520 88704
rect 4456 88644 4460 88700
rect 4460 88644 4516 88700
rect 4516 88644 4520 88700
rect 4456 88640 4520 88644
rect 34936 88700 35000 88704
rect 34936 88644 34940 88700
rect 34940 88644 34996 88700
rect 34996 88644 35000 88700
rect 34936 88640 35000 88644
rect 35016 88700 35080 88704
rect 35016 88644 35020 88700
rect 35020 88644 35076 88700
rect 35076 88644 35080 88700
rect 35016 88640 35080 88644
rect 35096 88700 35160 88704
rect 35096 88644 35100 88700
rect 35100 88644 35156 88700
rect 35156 88644 35160 88700
rect 35096 88640 35160 88644
rect 35176 88700 35240 88704
rect 35176 88644 35180 88700
rect 35180 88644 35236 88700
rect 35236 88644 35240 88700
rect 35176 88640 35240 88644
rect 65656 88700 65720 88704
rect 65656 88644 65660 88700
rect 65660 88644 65716 88700
rect 65716 88644 65720 88700
rect 65656 88640 65720 88644
rect 65736 88700 65800 88704
rect 65736 88644 65740 88700
rect 65740 88644 65796 88700
rect 65796 88644 65800 88700
rect 65736 88640 65800 88644
rect 65816 88700 65880 88704
rect 65816 88644 65820 88700
rect 65820 88644 65876 88700
rect 65876 88644 65880 88700
rect 65816 88640 65880 88644
rect 65896 88700 65960 88704
rect 65896 88644 65900 88700
rect 65900 88644 65956 88700
rect 65956 88644 65960 88700
rect 65896 88640 65960 88644
rect 96376 88700 96440 88704
rect 96376 88644 96380 88700
rect 96380 88644 96436 88700
rect 96436 88644 96440 88700
rect 96376 88640 96440 88644
rect 96456 88700 96520 88704
rect 96456 88644 96460 88700
rect 96460 88644 96516 88700
rect 96516 88644 96520 88700
rect 96456 88640 96520 88644
rect 96536 88700 96600 88704
rect 96536 88644 96540 88700
rect 96540 88644 96596 88700
rect 96596 88644 96600 88700
rect 96536 88640 96600 88644
rect 96616 88700 96680 88704
rect 96616 88644 96620 88700
rect 96620 88644 96676 88700
rect 96676 88644 96680 88700
rect 96616 88640 96680 88644
rect 4876 88156 4940 88160
rect 4876 88100 4880 88156
rect 4880 88100 4936 88156
rect 4936 88100 4940 88156
rect 4876 88096 4940 88100
rect 4956 88156 5020 88160
rect 4956 88100 4960 88156
rect 4960 88100 5016 88156
rect 5016 88100 5020 88156
rect 4956 88096 5020 88100
rect 5036 88156 5100 88160
rect 5036 88100 5040 88156
rect 5040 88100 5096 88156
rect 5096 88100 5100 88156
rect 5036 88096 5100 88100
rect 5116 88156 5180 88160
rect 5116 88100 5120 88156
rect 5120 88100 5176 88156
rect 5176 88100 5180 88156
rect 5116 88096 5180 88100
rect 35596 88156 35660 88160
rect 35596 88100 35600 88156
rect 35600 88100 35656 88156
rect 35656 88100 35660 88156
rect 35596 88096 35660 88100
rect 35676 88156 35740 88160
rect 35676 88100 35680 88156
rect 35680 88100 35736 88156
rect 35736 88100 35740 88156
rect 35676 88096 35740 88100
rect 35756 88156 35820 88160
rect 35756 88100 35760 88156
rect 35760 88100 35816 88156
rect 35816 88100 35820 88156
rect 35756 88096 35820 88100
rect 35836 88156 35900 88160
rect 35836 88100 35840 88156
rect 35840 88100 35896 88156
rect 35896 88100 35900 88156
rect 35836 88096 35900 88100
rect 66316 88156 66380 88160
rect 66316 88100 66320 88156
rect 66320 88100 66376 88156
rect 66376 88100 66380 88156
rect 66316 88096 66380 88100
rect 66396 88156 66460 88160
rect 66396 88100 66400 88156
rect 66400 88100 66456 88156
rect 66456 88100 66460 88156
rect 66396 88096 66460 88100
rect 66476 88156 66540 88160
rect 66476 88100 66480 88156
rect 66480 88100 66536 88156
rect 66536 88100 66540 88156
rect 66476 88096 66540 88100
rect 66556 88156 66620 88160
rect 66556 88100 66560 88156
rect 66560 88100 66616 88156
rect 66616 88100 66620 88156
rect 66556 88096 66620 88100
rect 97036 88156 97100 88160
rect 97036 88100 97040 88156
rect 97040 88100 97096 88156
rect 97096 88100 97100 88156
rect 97036 88096 97100 88100
rect 97116 88156 97180 88160
rect 97116 88100 97120 88156
rect 97120 88100 97176 88156
rect 97176 88100 97180 88156
rect 97116 88096 97180 88100
rect 97196 88156 97260 88160
rect 97196 88100 97200 88156
rect 97200 88100 97256 88156
rect 97256 88100 97260 88156
rect 97196 88096 97260 88100
rect 97276 88156 97340 88160
rect 97276 88100 97280 88156
rect 97280 88100 97336 88156
rect 97336 88100 97340 88156
rect 97276 88096 97340 88100
rect 4216 87612 4280 87616
rect 4216 87556 4220 87612
rect 4220 87556 4276 87612
rect 4276 87556 4280 87612
rect 4216 87552 4280 87556
rect 4296 87612 4360 87616
rect 4296 87556 4300 87612
rect 4300 87556 4356 87612
rect 4356 87556 4360 87612
rect 4296 87552 4360 87556
rect 4376 87612 4440 87616
rect 4376 87556 4380 87612
rect 4380 87556 4436 87612
rect 4436 87556 4440 87612
rect 4376 87552 4440 87556
rect 4456 87612 4520 87616
rect 4456 87556 4460 87612
rect 4460 87556 4516 87612
rect 4516 87556 4520 87612
rect 4456 87552 4520 87556
rect 34936 87612 35000 87616
rect 34936 87556 34940 87612
rect 34940 87556 34996 87612
rect 34996 87556 35000 87612
rect 34936 87552 35000 87556
rect 35016 87612 35080 87616
rect 35016 87556 35020 87612
rect 35020 87556 35076 87612
rect 35076 87556 35080 87612
rect 35016 87552 35080 87556
rect 35096 87612 35160 87616
rect 35096 87556 35100 87612
rect 35100 87556 35156 87612
rect 35156 87556 35160 87612
rect 35096 87552 35160 87556
rect 35176 87612 35240 87616
rect 35176 87556 35180 87612
rect 35180 87556 35236 87612
rect 35236 87556 35240 87612
rect 35176 87552 35240 87556
rect 65656 87612 65720 87616
rect 65656 87556 65660 87612
rect 65660 87556 65716 87612
rect 65716 87556 65720 87612
rect 65656 87552 65720 87556
rect 65736 87612 65800 87616
rect 65736 87556 65740 87612
rect 65740 87556 65796 87612
rect 65796 87556 65800 87612
rect 65736 87552 65800 87556
rect 65816 87612 65880 87616
rect 65816 87556 65820 87612
rect 65820 87556 65876 87612
rect 65876 87556 65880 87612
rect 65816 87552 65880 87556
rect 65896 87612 65960 87616
rect 65896 87556 65900 87612
rect 65900 87556 65956 87612
rect 65956 87556 65960 87612
rect 65896 87552 65960 87556
rect 96376 87612 96440 87616
rect 96376 87556 96380 87612
rect 96380 87556 96436 87612
rect 96436 87556 96440 87612
rect 96376 87552 96440 87556
rect 96456 87612 96520 87616
rect 96456 87556 96460 87612
rect 96460 87556 96516 87612
rect 96516 87556 96520 87612
rect 96456 87552 96520 87556
rect 96536 87612 96600 87616
rect 96536 87556 96540 87612
rect 96540 87556 96596 87612
rect 96596 87556 96600 87612
rect 96536 87552 96600 87556
rect 96616 87612 96680 87616
rect 96616 87556 96620 87612
rect 96620 87556 96676 87612
rect 96676 87556 96680 87612
rect 96616 87552 96680 87556
rect 4876 87068 4940 87072
rect 4876 87012 4880 87068
rect 4880 87012 4936 87068
rect 4936 87012 4940 87068
rect 4876 87008 4940 87012
rect 4956 87068 5020 87072
rect 4956 87012 4960 87068
rect 4960 87012 5016 87068
rect 5016 87012 5020 87068
rect 4956 87008 5020 87012
rect 5036 87068 5100 87072
rect 5036 87012 5040 87068
rect 5040 87012 5096 87068
rect 5096 87012 5100 87068
rect 5036 87008 5100 87012
rect 5116 87068 5180 87072
rect 5116 87012 5120 87068
rect 5120 87012 5176 87068
rect 5176 87012 5180 87068
rect 5116 87008 5180 87012
rect 35596 87068 35660 87072
rect 35596 87012 35600 87068
rect 35600 87012 35656 87068
rect 35656 87012 35660 87068
rect 35596 87008 35660 87012
rect 35676 87068 35740 87072
rect 35676 87012 35680 87068
rect 35680 87012 35736 87068
rect 35736 87012 35740 87068
rect 35676 87008 35740 87012
rect 35756 87068 35820 87072
rect 35756 87012 35760 87068
rect 35760 87012 35816 87068
rect 35816 87012 35820 87068
rect 35756 87008 35820 87012
rect 35836 87068 35900 87072
rect 35836 87012 35840 87068
rect 35840 87012 35896 87068
rect 35896 87012 35900 87068
rect 35836 87008 35900 87012
rect 66316 87068 66380 87072
rect 66316 87012 66320 87068
rect 66320 87012 66376 87068
rect 66376 87012 66380 87068
rect 66316 87008 66380 87012
rect 66396 87068 66460 87072
rect 66396 87012 66400 87068
rect 66400 87012 66456 87068
rect 66456 87012 66460 87068
rect 66396 87008 66460 87012
rect 66476 87068 66540 87072
rect 66476 87012 66480 87068
rect 66480 87012 66536 87068
rect 66536 87012 66540 87068
rect 66476 87008 66540 87012
rect 66556 87068 66620 87072
rect 66556 87012 66560 87068
rect 66560 87012 66616 87068
rect 66616 87012 66620 87068
rect 66556 87008 66620 87012
rect 97036 87068 97100 87072
rect 97036 87012 97040 87068
rect 97040 87012 97096 87068
rect 97096 87012 97100 87068
rect 97036 87008 97100 87012
rect 97116 87068 97180 87072
rect 97116 87012 97120 87068
rect 97120 87012 97176 87068
rect 97176 87012 97180 87068
rect 97116 87008 97180 87012
rect 97196 87068 97260 87072
rect 97196 87012 97200 87068
rect 97200 87012 97256 87068
rect 97256 87012 97260 87068
rect 97196 87008 97260 87012
rect 97276 87068 97340 87072
rect 97276 87012 97280 87068
rect 97280 87012 97336 87068
rect 97336 87012 97340 87068
rect 97276 87008 97340 87012
rect 4216 86524 4280 86528
rect 4216 86468 4220 86524
rect 4220 86468 4276 86524
rect 4276 86468 4280 86524
rect 4216 86464 4280 86468
rect 4296 86524 4360 86528
rect 4296 86468 4300 86524
rect 4300 86468 4356 86524
rect 4356 86468 4360 86524
rect 4296 86464 4360 86468
rect 4376 86524 4440 86528
rect 4376 86468 4380 86524
rect 4380 86468 4436 86524
rect 4436 86468 4440 86524
rect 4376 86464 4440 86468
rect 4456 86524 4520 86528
rect 4456 86468 4460 86524
rect 4460 86468 4516 86524
rect 4516 86468 4520 86524
rect 4456 86464 4520 86468
rect 34936 86524 35000 86528
rect 34936 86468 34940 86524
rect 34940 86468 34996 86524
rect 34996 86468 35000 86524
rect 34936 86464 35000 86468
rect 35016 86524 35080 86528
rect 35016 86468 35020 86524
rect 35020 86468 35076 86524
rect 35076 86468 35080 86524
rect 35016 86464 35080 86468
rect 35096 86524 35160 86528
rect 35096 86468 35100 86524
rect 35100 86468 35156 86524
rect 35156 86468 35160 86524
rect 35096 86464 35160 86468
rect 35176 86524 35240 86528
rect 35176 86468 35180 86524
rect 35180 86468 35236 86524
rect 35236 86468 35240 86524
rect 35176 86464 35240 86468
rect 65656 86524 65720 86528
rect 65656 86468 65660 86524
rect 65660 86468 65716 86524
rect 65716 86468 65720 86524
rect 65656 86464 65720 86468
rect 65736 86524 65800 86528
rect 65736 86468 65740 86524
rect 65740 86468 65796 86524
rect 65796 86468 65800 86524
rect 65736 86464 65800 86468
rect 65816 86524 65880 86528
rect 65816 86468 65820 86524
rect 65820 86468 65876 86524
rect 65876 86468 65880 86524
rect 65816 86464 65880 86468
rect 65896 86524 65960 86528
rect 65896 86468 65900 86524
rect 65900 86468 65956 86524
rect 65956 86468 65960 86524
rect 65896 86464 65960 86468
rect 96376 86524 96440 86528
rect 96376 86468 96380 86524
rect 96380 86468 96436 86524
rect 96436 86468 96440 86524
rect 96376 86464 96440 86468
rect 96456 86524 96520 86528
rect 96456 86468 96460 86524
rect 96460 86468 96516 86524
rect 96516 86468 96520 86524
rect 96456 86464 96520 86468
rect 96536 86524 96600 86528
rect 96536 86468 96540 86524
rect 96540 86468 96596 86524
rect 96596 86468 96600 86524
rect 96536 86464 96600 86468
rect 96616 86524 96680 86528
rect 96616 86468 96620 86524
rect 96620 86468 96676 86524
rect 96676 86468 96680 86524
rect 96616 86464 96680 86468
rect 4876 85980 4940 85984
rect 4876 85924 4880 85980
rect 4880 85924 4936 85980
rect 4936 85924 4940 85980
rect 4876 85920 4940 85924
rect 4956 85980 5020 85984
rect 4956 85924 4960 85980
rect 4960 85924 5016 85980
rect 5016 85924 5020 85980
rect 4956 85920 5020 85924
rect 5036 85980 5100 85984
rect 5036 85924 5040 85980
rect 5040 85924 5096 85980
rect 5096 85924 5100 85980
rect 5036 85920 5100 85924
rect 5116 85980 5180 85984
rect 5116 85924 5120 85980
rect 5120 85924 5176 85980
rect 5176 85924 5180 85980
rect 5116 85920 5180 85924
rect 35596 85980 35660 85984
rect 35596 85924 35600 85980
rect 35600 85924 35656 85980
rect 35656 85924 35660 85980
rect 35596 85920 35660 85924
rect 35676 85980 35740 85984
rect 35676 85924 35680 85980
rect 35680 85924 35736 85980
rect 35736 85924 35740 85980
rect 35676 85920 35740 85924
rect 35756 85980 35820 85984
rect 35756 85924 35760 85980
rect 35760 85924 35816 85980
rect 35816 85924 35820 85980
rect 35756 85920 35820 85924
rect 35836 85980 35900 85984
rect 35836 85924 35840 85980
rect 35840 85924 35896 85980
rect 35896 85924 35900 85980
rect 35836 85920 35900 85924
rect 66316 85980 66380 85984
rect 66316 85924 66320 85980
rect 66320 85924 66376 85980
rect 66376 85924 66380 85980
rect 66316 85920 66380 85924
rect 66396 85980 66460 85984
rect 66396 85924 66400 85980
rect 66400 85924 66456 85980
rect 66456 85924 66460 85980
rect 66396 85920 66460 85924
rect 66476 85980 66540 85984
rect 66476 85924 66480 85980
rect 66480 85924 66536 85980
rect 66536 85924 66540 85980
rect 66476 85920 66540 85924
rect 66556 85980 66620 85984
rect 66556 85924 66560 85980
rect 66560 85924 66616 85980
rect 66616 85924 66620 85980
rect 66556 85920 66620 85924
rect 97036 85980 97100 85984
rect 97036 85924 97040 85980
rect 97040 85924 97096 85980
rect 97096 85924 97100 85980
rect 97036 85920 97100 85924
rect 97116 85980 97180 85984
rect 97116 85924 97120 85980
rect 97120 85924 97176 85980
rect 97176 85924 97180 85980
rect 97116 85920 97180 85924
rect 97196 85980 97260 85984
rect 97196 85924 97200 85980
rect 97200 85924 97256 85980
rect 97256 85924 97260 85980
rect 97196 85920 97260 85924
rect 97276 85980 97340 85984
rect 97276 85924 97280 85980
rect 97280 85924 97336 85980
rect 97336 85924 97340 85980
rect 97276 85920 97340 85924
rect 4216 85436 4280 85440
rect 4216 85380 4220 85436
rect 4220 85380 4276 85436
rect 4276 85380 4280 85436
rect 4216 85376 4280 85380
rect 4296 85436 4360 85440
rect 4296 85380 4300 85436
rect 4300 85380 4356 85436
rect 4356 85380 4360 85436
rect 4296 85376 4360 85380
rect 4376 85436 4440 85440
rect 4376 85380 4380 85436
rect 4380 85380 4436 85436
rect 4436 85380 4440 85436
rect 4376 85376 4440 85380
rect 4456 85436 4520 85440
rect 4456 85380 4460 85436
rect 4460 85380 4516 85436
rect 4516 85380 4520 85436
rect 4456 85376 4520 85380
rect 34936 85436 35000 85440
rect 34936 85380 34940 85436
rect 34940 85380 34996 85436
rect 34996 85380 35000 85436
rect 34936 85376 35000 85380
rect 35016 85436 35080 85440
rect 35016 85380 35020 85436
rect 35020 85380 35076 85436
rect 35076 85380 35080 85436
rect 35016 85376 35080 85380
rect 35096 85436 35160 85440
rect 35096 85380 35100 85436
rect 35100 85380 35156 85436
rect 35156 85380 35160 85436
rect 35096 85376 35160 85380
rect 35176 85436 35240 85440
rect 35176 85380 35180 85436
rect 35180 85380 35236 85436
rect 35236 85380 35240 85436
rect 35176 85376 35240 85380
rect 65656 85436 65720 85440
rect 65656 85380 65660 85436
rect 65660 85380 65716 85436
rect 65716 85380 65720 85436
rect 65656 85376 65720 85380
rect 65736 85436 65800 85440
rect 65736 85380 65740 85436
rect 65740 85380 65796 85436
rect 65796 85380 65800 85436
rect 65736 85376 65800 85380
rect 65816 85436 65880 85440
rect 65816 85380 65820 85436
rect 65820 85380 65876 85436
rect 65876 85380 65880 85436
rect 65816 85376 65880 85380
rect 65896 85436 65960 85440
rect 65896 85380 65900 85436
rect 65900 85380 65956 85436
rect 65956 85380 65960 85436
rect 65896 85376 65960 85380
rect 96376 85436 96440 85440
rect 96376 85380 96380 85436
rect 96380 85380 96436 85436
rect 96436 85380 96440 85436
rect 96376 85376 96440 85380
rect 96456 85436 96520 85440
rect 96456 85380 96460 85436
rect 96460 85380 96516 85436
rect 96516 85380 96520 85436
rect 96456 85376 96520 85380
rect 96536 85436 96600 85440
rect 96536 85380 96540 85436
rect 96540 85380 96596 85436
rect 96596 85380 96600 85436
rect 96536 85376 96600 85380
rect 96616 85436 96680 85440
rect 96616 85380 96620 85436
rect 96620 85380 96676 85436
rect 96676 85380 96680 85436
rect 96616 85376 96680 85380
rect 4876 84892 4940 84896
rect 4876 84836 4880 84892
rect 4880 84836 4936 84892
rect 4936 84836 4940 84892
rect 4876 84832 4940 84836
rect 4956 84892 5020 84896
rect 4956 84836 4960 84892
rect 4960 84836 5016 84892
rect 5016 84836 5020 84892
rect 4956 84832 5020 84836
rect 5036 84892 5100 84896
rect 5036 84836 5040 84892
rect 5040 84836 5096 84892
rect 5096 84836 5100 84892
rect 5036 84832 5100 84836
rect 5116 84892 5180 84896
rect 5116 84836 5120 84892
rect 5120 84836 5176 84892
rect 5176 84836 5180 84892
rect 5116 84832 5180 84836
rect 35596 84892 35660 84896
rect 35596 84836 35600 84892
rect 35600 84836 35656 84892
rect 35656 84836 35660 84892
rect 35596 84832 35660 84836
rect 35676 84892 35740 84896
rect 35676 84836 35680 84892
rect 35680 84836 35736 84892
rect 35736 84836 35740 84892
rect 35676 84832 35740 84836
rect 35756 84892 35820 84896
rect 35756 84836 35760 84892
rect 35760 84836 35816 84892
rect 35816 84836 35820 84892
rect 35756 84832 35820 84836
rect 35836 84892 35900 84896
rect 35836 84836 35840 84892
rect 35840 84836 35896 84892
rect 35896 84836 35900 84892
rect 35836 84832 35900 84836
rect 66316 84892 66380 84896
rect 66316 84836 66320 84892
rect 66320 84836 66376 84892
rect 66376 84836 66380 84892
rect 66316 84832 66380 84836
rect 66396 84892 66460 84896
rect 66396 84836 66400 84892
rect 66400 84836 66456 84892
rect 66456 84836 66460 84892
rect 66396 84832 66460 84836
rect 66476 84892 66540 84896
rect 66476 84836 66480 84892
rect 66480 84836 66536 84892
rect 66536 84836 66540 84892
rect 66476 84832 66540 84836
rect 66556 84892 66620 84896
rect 66556 84836 66560 84892
rect 66560 84836 66616 84892
rect 66616 84836 66620 84892
rect 66556 84832 66620 84836
rect 97036 84892 97100 84896
rect 97036 84836 97040 84892
rect 97040 84836 97096 84892
rect 97096 84836 97100 84892
rect 97036 84832 97100 84836
rect 97116 84892 97180 84896
rect 97116 84836 97120 84892
rect 97120 84836 97176 84892
rect 97176 84836 97180 84892
rect 97116 84832 97180 84836
rect 97196 84892 97260 84896
rect 97196 84836 97200 84892
rect 97200 84836 97256 84892
rect 97256 84836 97260 84892
rect 97196 84832 97260 84836
rect 97276 84892 97340 84896
rect 97276 84836 97280 84892
rect 97280 84836 97336 84892
rect 97336 84836 97340 84892
rect 97276 84832 97340 84836
rect 4216 84348 4280 84352
rect 4216 84292 4220 84348
rect 4220 84292 4276 84348
rect 4276 84292 4280 84348
rect 4216 84288 4280 84292
rect 4296 84348 4360 84352
rect 4296 84292 4300 84348
rect 4300 84292 4356 84348
rect 4356 84292 4360 84348
rect 4296 84288 4360 84292
rect 4376 84348 4440 84352
rect 4376 84292 4380 84348
rect 4380 84292 4436 84348
rect 4436 84292 4440 84348
rect 4376 84288 4440 84292
rect 4456 84348 4520 84352
rect 4456 84292 4460 84348
rect 4460 84292 4516 84348
rect 4516 84292 4520 84348
rect 4456 84288 4520 84292
rect 34936 84348 35000 84352
rect 34936 84292 34940 84348
rect 34940 84292 34996 84348
rect 34996 84292 35000 84348
rect 34936 84288 35000 84292
rect 35016 84348 35080 84352
rect 35016 84292 35020 84348
rect 35020 84292 35076 84348
rect 35076 84292 35080 84348
rect 35016 84288 35080 84292
rect 35096 84348 35160 84352
rect 35096 84292 35100 84348
rect 35100 84292 35156 84348
rect 35156 84292 35160 84348
rect 35096 84288 35160 84292
rect 35176 84348 35240 84352
rect 35176 84292 35180 84348
rect 35180 84292 35236 84348
rect 35236 84292 35240 84348
rect 35176 84288 35240 84292
rect 65656 84348 65720 84352
rect 65656 84292 65660 84348
rect 65660 84292 65716 84348
rect 65716 84292 65720 84348
rect 65656 84288 65720 84292
rect 65736 84348 65800 84352
rect 65736 84292 65740 84348
rect 65740 84292 65796 84348
rect 65796 84292 65800 84348
rect 65736 84288 65800 84292
rect 65816 84348 65880 84352
rect 65816 84292 65820 84348
rect 65820 84292 65876 84348
rect 65876 84292 65880 84348
rect 65816 84288 65880 84292
rect 65896 84348 65960 84352
rect 65896 84292 65900 84348
rect 65900 84292 65956 84348
rect 65956 84292 65960 84348
rect 65896 84288 65960 84292
rect 96376 84348 96440 84352
rect 96376 84292 96380 84348
rect 96380 84292 96436 84348
rect 96436 84292 96440 84348
rect 96376 84288 96440 84292
rect 96456 84348 96520 84352
rect 96456 84292 96460 84348
rect 96460 84292 96516 84348
rect 96516 84292 96520 84348
rect 96456 84288 96520 84292
rect 96536 84348 96600 84352
rect 96536 84292 96540 84348
rect 96540 84292 96596 84348
rect 96596 84292 96600 84348
rect 96536 84288 96600 84292
rect 96616 84348 96680 84352
rect 96616 84292 96620 84348
rect 96620 84292 96676 84348
rect 96676 84292 96680 84348
rect 96616 84288 96680 84292
rect 4876 83804 4940 83808
rect 4876 83748 4880 83804
rect 4880 83748 4936 83804
rect 4936 83748 4940 83804
rect 4876 83744 4940 83748
rect 4956 83804 5020 83808
rect 4956 83748 4960 83804
rect 4960 83748 5016 83804
rect 5016 83748 5020 83804
rect 4956 83744 5020 83748
rect 5036 83804 5100 83808
rect 5036 83748 5040 83804
rect 5040 83748 5096 83804
rect 5096 83748 5100 83804
rect 5036 83744 5100 83748
rect 5116 83804 5180 83808
rect 5116 83748 5120 83804
rect 5120 83748 5176 83804
rect 5176 83748 5180 83804
rect 5116 83744 5180 83748
rect 35596 83804 35660 83808
rect 35596 83748 35600 83804
rect 35600 83748 35656 83804
rect 35656 83748 35660 83804
rect 35596 83744 35660 83748
rect 35676 83804 35740 83808
rect 35676 83748 35680 83804
rect 35680 83748 35736 83804
rect 35736 83748 35740 83804
rect 35676 83744 35740 83748
rect 35756 83804 35820 83808
rect 35756 83748 35760 83804
rect 35760 83748 35816 83804
rect 35816 83748 35820 83804
rect 35756 83744 35820 83748
rect 35836 83804 35900 83808
rect 35836 83748 35840 83804
rect 35840 83748 35896 83804
rect 35896 83748 35900 83804
rect 35836 83744 35900 83748
rect 66316 83804 66380 83808
rect 66316 83748 66320 83804
rect 66320 83748 66376 83804
rect 66376 83748 66380 83804
rect 66316 83744 66380 83748
rect 66396 83804 66460 83808
rect 66396 83748 66400 83804
rect 66400 83748 66456 83804
rect 66456 83748 66460 83804
rect 66396 83744 66460 83748
rect 66476 83804 66540 83808
rect 66476 83748 66480 83804
rect 66480 83748 66536 83804
rect 66536 83748 66540 83804
rect 66476 83744 66540 83748
rect 66556 83804 66620 83808
rect 66556 83748 66560 83804
rect 66560 83748 66616 83804
rect 66616 83748 66620 83804
rect 66556 83744 66620 83748
rect 97036 83804 97100 83808
rect 97036 83748 97040 83804
rect 97040 83748 97096 83804
rect 97096 83748 97100 83804
rect 97036 83744 97100 83748
rect 97116 83804 97180 83808
rect 97116 83748 97120 83804
rect 97120 83748 97176 83804
rect 97176 83748 97180 83804
rect 97116 83744 97180 83748
rect 97196 83804 97260 83808
rect 97196 83748 97200 83804
rect 97200 83748 97256 83804
rect 97256 83748 97260 83804
rect 97196 83744 97260 83748
rect 97276 83804 97340 83808
rect 97276 83748 97280 83804
rect 97280 83748 97336 83804
rect 97336 83748 97340 83804
rect 97276 83744 97340 83748
rect 4216 83260 4280 83264
rect 4216 83204 4220 83260
rect 4220 83204 4276 83260
rect 4276 83204 4280 83260
rect 4216 83200 4280 83204
rect 4296 83260 4360 83264
rect 4296 83204 4300 83260
rect 4300 83204 4356 83260
rect 4356 83204 4360 83260
rect 4296 83200 4360 83204
rect 4376 83260 4440 83264
rect 4376 83204 4380 83260
rect 4380 83204 4436 83260
rect 4436 83204 4440 83260
rect 4376 83200 4440 83204
rect 4456 83260 4520 83264
rect 4456 83204 4460 83260
rect 4460 83204 4516 83260
rect 4516 83204 4520 83260
rect 4456 83200 4520 83204
rect 34936 83260 35000 83264
rect 34936 83204 34940 83260
rect 34940 83204 34996 83260
rect 34996 83204 35000 83260
rect 34936 83200 35000 83204
rect 35016 83260 35080 83264
rect 35016 83204 35020 83260
rect 35020 83204 35076 83260
rect 35076 83204 35080 83260
rect 35016 83200 35080 83204
rect 35096 83260 35160 83264
rect 35096 83204 35100 83260
rect 35100 83204 35156 83260
rect 35156 83204 35160 83260
rect 35096 83200 35160 83204
rect 35176 83260 35240 83264
rect 35176 83204 35180 83260
rect 35180 83204 35236 83260
rect 35236 83204 35240 83260
rect 35176 83200 35240 83204
rect 65656 83260 65720 83264
rect 65656 83204 65660 83260
rect 65660 83204 65716 83260
rect 65716 83204 65720 83260
rect 65656 83200 65720 83204
rect 65736 83260 65800 83264
rect 65736 83204 65740 83260
rect 65740 83204 65796 83260
rect 65796 83204 65800 83260
rect 65736 83200 65800 83204
rect 65816 83260 65880 83264
rect 65816 83204 65820 83260
rect 65820 83204 65876 83260
rect 65876 83204 65880 83260
rect 65816 83200 65880 83204
rect 65896 83260 65960 83264
rect 65896 83204 65900 83260
rect 65900 83204 65956 83260
rect 65956 83204 65960 83260
rect 65896 83200 65960 83204
rect 96376 83260 96440 83264
rect 96376 83204 96380 83260
rect 96380 83204 96436 83260
rect 96436 83204 96440 83260
rect 96376 83200 96440 83204
rect 96456 83260 96520 83264
rect 96456 83204 96460 83260
rect 96460 83204 96516 83260
rect 96516 83204 96520 83260
rect 96456 83200 96520 83204
rect 96536 83260 96600 83264
rect 96536 83204 96540 83260
rect 96540 83204 96596 83260
rect 96596 83204 96600 83260
rect 96536 83200 96600 83204
rect 96616 83260 96680 83264
rect 96616 83204 96620 83260
rect 96620 83204 96676 83260
rect 96676 83204 96680 83260
rect 96616 83200 96680 83204
rect 4876 82716 4940 82720
rect 4876 82660 4880 82716
rect 4880 82660 4936 82716
rect 4936 82660 4940 82716
rect 4876 82656 4940 82660
rect 4956 82716 5020 82720
rect 4956 82660 4960 82716
rect 4960 82660 5016 82716
rect 5016 82660 5020 82716
rect 4956 82656 5020 82660
rect 5036 82716 5100 82720
rect 5036 82660 5040 82716
rect 5040 82660 5096 82716
rect 5096 82660 5100 82716
rect 5036 82656 5100 82660
rect 5116 82716 5180 82720
rect 5116 82660 5120 82716
rect 5120 82660 5176 82716
rect 5176 82660 5180 82716
rect 5116 82656 5180 82660
rect 35596 82716 35660 82720
rect 35596 82660 35600 82716
rect 35600 82660 35656 82716
rect 35656 82660 35660 82716
rect 35596 82656 35660 82660
rect 35676 82716 35740 82720
rect 35676 82660 35680 82716
rect 35680 82660 35736 82716
rect 35736 82660 35740 82716
rect 35676 82656 35740 82660
rect 35756 82716 35820 82720
rect 35756 82660 35760 82716
rect 35760 82660 35816 82716
rect 35816 82660 35820 82716
rect 35756 82656 35820 82660
rect 35836 82716 35900 82720
rect 35836 82660 35840 82716
rect 35840 82660 35896 82716
rect 35896 82660 35900 82716
rect 35836 82656 35900 82660
rect 66316 82716 66380 82720
rect 66316 82660 66320 82716
rect 66320 82660 66376 82716
rect 66376 82660 66380 82716
rect 66316 82656 66380 82660
rect 66396 82716 66460 82720
rect 66396 82660 66400 82716
rect 66400 82660 66456 82716
rect 66456 82660 66460 82716
rect 66396 82656 66460 82660
rect 66476 82716 66540 82720
rect 66476 82660 66480 82716
rect 66480 82660 66536 82716
rect 66536 82660 66540 82716
rect 66476 82656 66540 82660
rect 66556 82716 66620 82720
rect 66556 82660 66560 82716
rect 66560 82660 66616 82716
rect 66616 82660 66620 82716
rect 66556 82656 66620 82660
rect 97036 82716 97100 82720
rect 97036 82660 97040 82716
rect 97040 82660 97096 82716
rect 97096 82660 97100 82716
rect 97036 82656 97100 82660
rect 97116 82716 97180 82720
rect 97116 82660 97120 82716
rect 97120 82660 97176 82716
rect 97176 82660 97180 82716
rect 97116 82656 97180 82660
rect 97196 82716 97260 82720
rect 97196 82660 97200 82716
rect 97200 82660 97256 82716
rect 97256 82660 97260 82716
rect 97196 82656 97260 82660
rect 97276 82716 97340 82720
rect 97276 82660 97280 82716
rect 97280 82660 97336 82716
rect 97336 82660 97340 82716
rect 97276 82656 97340 82660
rect 4216 82172 4280 82176
rect 4216 82116 4220 82172
rect 4220 82116 4276 82172
rect 4276 82116 4280 82172
rect 4216 82112 4280 82116
rect 4296 82172 4360 82176
rect 4296 82116 4300 82172
rect 4300 82116 4356 82172
rect 4356 82116 4360 82172
rect 4296 82112 4360 82116
rect 4376 82172 4440 82176
rect 4376 82116 4380 82172
rect 4380 82116 4436 82172
rect 4436 82116 4440 82172
rect 4376 82112 4440 82116
rect 4456 82172 4520 82176
rect 4456 82116 4460 82172
rect 4460 82116 4516 82172
rect 4516 82116 4520 82172
rect 4456 82112 4520 82116
rect 34936 82172 35000 82176
rect 34936 82116 34940 82172
rect 34940 82116 34996 82172
rect 34996 82116 35000 82172
rect 34936 82112 35000 82116
rect 35016 82172 35080 82176
rect 35016 82116 35020 82172
rect 35020 82116 35076 82172
rect 35076 82116 35080 82172
rect 35016 82112 35080 82116
rect 35096 82172 35160 82176
rect 35096 82116 35100 82172
rect 35100 82116 35156 82172
rect 35156 82116 35160 82172
rect 35096 82112 35160 82116
rect 35176 82172 35240 82176
rect 35176 82116 35180 82172
rect 35180 82116 35236 82172
rect 35236 82116 35240 82172
rect 35176 82112 35240 82116
rect 65656 82172 65720 82176
rect 65656 82116 65660 82172
rect 65660 82116 65716 82172
rect 65716 82116 65720 82172
rect 65656 82112 65720 82116
rect 65736 82172 65800 82176
rect 65736 82116 65740 82172
rect 65740 82116 65796 82172
rect 65796 82116 65800 82172
rect 65736 82112 65800 82116
rect 65816 82172 65880 82176
rect 65816 82116 65820 82172
rect 65820 82116 65876 82172
rect 65876 82116 65880 82172
rect 65816 82112 65880 82116
rect 65896 82172 65960 82176
rect 65896 82116 65900 82172
rect 65900 82116 65956 82172
rect 65956 82116 65960 82172
rect 65896 82112 65960 82116
rect 96376 82172 96440 82176
rect 96376 82116 96380 82172
rect 96380 82116 96436 82172
rect 96436 82116 96440 82172
rect 96376 82112 96440 82116
rect 96456 82172 96520 82176
rect 96456 82116 96460 82172
rect 96460 82116 96516 82172
rect 96516 82116 96520 82172
rect 96456 82112 96520 82116
rect 96536 82172 96600 82176
rect 96536 82116 96540 82172
rect 96540 82116 96596 82172
rect 96596 82116 96600 82172
rect 96536 82112 96600 82116
rect 96616 82172 96680 82176
rect 96616 82116 96620 82172
rect 96620 82116 96676 82172
rect 96676 82116 96680 82172
rect 96616 82112 96680 82116
rect 4876 81628 4940 81632
rect 4876 81572 4880 81628
rect 4880 81572 4936 81628
rect 4936 81572 4940 81628
rect 4876 81568 4940 81572
rect 4956 81628 5020 81632
rect 4956 81572 4960 81628
rect 4960 81572 5016 81628
rect 5016 81572 5020 81628
rect 4956 81568 5020 81572
rect 5036 81628 5100 81632
rect 5036 81572 5040 81628
rect 5040 81572 5096 81628
rect 5096 81572 5100 81628
rect 5036 81568 5100 81572
rect 5116 81628 5180 81632
rect 5116 81572 5120 81628
rect 5120 81572 5176 81628
rect 5176 81572 5180 81628
rect 5116 81568 5180 81572
rect 35596 81628 35660 81632
rect 35596 81572 35600 81628
rect 35600 81572 35656 81628
rect 35656 81572 35660 81628
rect 35596 81568 35660 81572
rect 35676 81628 35740 81632
rect 35676 81572 35680 81628
rect 35680 81572 35736 81628
rect 35736 81572 35740 81628
rect 35676 81568 35740 81572
rect 35756 81628 35820 81632
rect 35756 81572 35760 81628
rect 35760 81572 35816 81628
rect 35816 81572 35820 81628
rect 35756 81568 35820 81572
rect 35836 81628 35900 81632
rect 35836 81572 35840 81628
rect 35840 81572 35896 81628
rect 35896 81572 35900 81628
rect 35836 81568 35900 81572
rect 66316 81628 66380 81632
rect 66316 81572 66320 81628
rect 66320 81572 66376 81628
rect 66376 81572 66380 81628
rect 66316 81568 66380 81572
rect 66396 81628 66460 81632
rect 66396 81572 66400 81628
rect 66400 81572 66456 81628
rect 66456 81572 66460 81628
rect 66396 81568 66460 81572
rect 66476 81628 66540 81632
rect 66476 81572 66480 81628
rect 66480 81572 66536 81628
rect 66536 81572 66540 81628
rect 66476 81568 66540 81572
rect 66556 81628 66620 81632
rect 66556 81572 66560 81628
rect 66560 81572 66616 81628
rect 66616 81572 66620 81628
rect 66556 81568 66620 81572
rect 97036 81628 97100 81632
rect 97036 81572 97040 81628
rect 97040 81572 97096 81628
rect 97096 81572 97100 81628
rect 97036 81568 97100 81572
rect 97116 81628 97180 81632
rect 97116 81572 97120 81628
rect 97120 81572 97176 81628
rect 97176 81572 97180 81628
rect 97116 81568 97180 81572
rect 97196 81628 97260 81632
rect 97196 81572 97200 81628
rect 97200 81572 97256 81628
rect 97256 81572 97260 81628
rect 97196 81568 97260 81572
rect 97276 81628 97340 81632
rect 97276 81572 97280 81628
rect 97280 81572 97336 81628
rect 97336 81572 97340 81628
rect 97276 81568 97340 81572
rect 4216 81084 4280 81088
rect 4216 81028 4220 81084
rect 4220 81028 4276 81084
rect 4276 81028 4280 81084
rect 4216 81024 4280 81028
rect 4296 81084 4360 81088
rect 4296 81028 4300 81084
rect 4300 81028 4356 81084
rect 4356 81028 4360 81084
rect 4296 81024 4360 81028
rect 4376 81084 4440 81088
rect 4376 81028 4380 81084
rect 4380 81028 4436 81084
rect 4436 81028 4440 81084
rect 4376 81024 4440 81028
rect 4456 81084 4520 81088
rect 4456 81028 4460 81084
rect 4460 81028 4516 81084
rect 4516 81028 4520 81084
rect 4456 81024 4520 81028
rect 34936 81084 35000 81088
rect 34936 81028 34940 81084
rect 34940 81028 34996 81084
rect 34996 81028 35000 81084
rect 34936 81024 35000 81028
rect 35016 81084 35080 81088
rect 35016 81028 35020 81084
rect 35020 81028 35076 81084
rect 35076 81028 35080 81084
rect 35016 81024 35080 81028
rect 35096 81084 35160 81088
rect 35096 81028 35100 81084
rect 35100 81028 35156 81084
rect 35156 81028 35160 81084
rect 35096 81024 35160 81028
rect 35176 81084 35240 81088
rect 35176 81028 35180 81084
rect 35180 81028 35236 81084
rect 35236 81028 35240 81084
rect 35176 81024 35240 81028
rect 65656 81084 65720 81088
rect 65656 81028 65660 81084
rect 65660 81028 65716 81084
rect 65716 81028 65720 81084
rect 65656 81024 65720 81028
rect 65736 81084 65800 81088
rect 65736 81028 65740 81084
rect 65740 81028 65796 81084
rect 65796 81028 65800 81084
rect 65736 81024 65800 81028
rect 65816 81084 65880 81088
rect 65816 81028 65820 81084
rect 65820 81028 65876 81084
rect 65876 81028 65880 81084
rect 65816 81024 65880 81028
rect 65896 81084 65960 81088
rect 65896 81028 65900 81084
rect 65900 81028 65956 81084
rect 65956 81028 65960 81084
rect 65896 81024 65960 81028
rect 96376 81084 96440 81088
rect 96376 81028 96380 81084
rect 96380 81028 96436 81084
rect 96436 81028 96440 81084
rect 96376 81024 96440 81028
rect 96456 81084 96520 81088
rect 96456 81028 96460 81084
rect 96460 81028 96516 81084
rect 96516 81028 96520 81084
rect 96456 81024 96520 81028
rect 96536 81084 96600 81088
rect 96536 81028 96540 81084
rect 96540 81028 96596 81084
rect 96596 81028 96600 81084
rect 96536 81024 96600 81028
rect 96616 81084 96680 81088
rect 96616 81028 96620 81084
rect 96620 81028 96676 81084
rect 96676 81028 96680 81084
rect 96616 81024 96680 81028
rect 4876 80540 4940 80544
rect 4876 80484 4880 80540
rect 4880 80484 4936 80540
rect 4936 80484 4940 80540
rect 4876 80480 4940 80484
rect 4956 80540 5020 80544
rect 4956 80484 4960 80540
rect 4960 80484 5016 80540
rect 5016 80484 5020 80540
rect 4956 80480 5020 80484
rect 5036 80540 5100 80544
rect 5036 80484 5040 80540
rect 5040 80484 5096 80540
rect 5096 80484 5100 80540
rect 5036 80480 5100 80484
rect 5116 80540 5180 80544
rect 5116 80484 5120 80540
rect 5120 80484 5176 80540
rect 5176 80484 5180 80540
rect 5116 80480 5180 80484
rect 35596 80540 35660 80544
rect 35596 80484 35600 80540
rect 35600 80484 35656 80540
rect 35656 80484 35660 80540
rect 35596 80480 35660 80484
rect 35676 80540 35740 80544
rect 35676 80484 35680 80540
rect 35680 80484 35736 80540
rect 35736 80484 35740 80540
rect 35676 80480 35740 80484
rect 35756 80540 35820 80544
rect 35756 80484 35760 80540
rect 35760 80484 35816 80540
rect 35816 80484 35820 80540
rect 35756 80480 35820 80484
rect 35836 80540 35900 80544
rect 35836 80484 35840 80540
rect 35840 80484 35896 80540
rect 35896 80484 35900 80540
rect 35836 80480 35900 80484
rect 66316 80540 66380 80544
rect 66316 80484 66320 80540
rect 66320 80484 66376 80540
rect 66376 80484 66380 80540
rect 66316 80480 66380 80484
rect 66396 80540 66460 80544
rect 66396 80484 66400 80540
rect 66400 80484 66456 80540
rect 66456 80484 66460 80540
rect 66396 80480 66460 80484
rect 66476 80540 66540 80544
rect 66476 80484 66480 80540
rect 66480 80484 66536 80540
rect 66536 80484 66540 80540
rect 66476 80480 66540 80484
rect 66556 80540 66620 80544
rect 66556 80484 66560 80540
rect 66560 80484 66616 80540
rect 66616 80484 66620 80540
rect 66556 80480 66620 80484
rect 97036 80540 97100 80544
rect 97036 80484 97040 80540
rect 97040 80484 97096 80540
rect 97096 80484 97100 80540
rect 97036 80480 97100 80484
rect 97116 80540 97180 80544
rect 97116 80484 97120 80540
rect 97120 80484 97176 80540
rect 97176 80484 97180 80540
rect 97116 80480 97180 80484
rect 97196 80540 97260 80544
rect 97196 80484 97200 80540
rect 97200 80484 97256 80540
rect 97256 80484 97260 80540
rect 97196 80480 97260 80484
rect 97276 80540 97340 80544
rect 97276 80484 97280 80540
rect 97280 80484 97336 80540
rect 97336 80484 97340 80540
rect 97276 80480 97340 80484
rect 4216 79996 4280 80000
rect 4216 79940 4220 79996
rect 4220 79940 4276 79996
rect 4276 79940 4280 79996
rect 4216 79936 4280 79940
rect 4296 79996 4360 80000
rect 4296 79940 4300 79996
rect 4300 79940 4356 79996
rect 4356 79940 4360 79996
rect 4296 79936 4360 79940
rect 4376 79996 4440 80000
rect 4376 79940 4380 79996
rect 4380 79940 4436 79996
rect 4436 79940 4440 79996
rect 4376 79936 4440 79940
rect 4456 79996 4520 80000
rect 4456 79940 4460 79996
rect 4460 79940 4516 79996
rect 4516 79940 4520 79996
rect 4456 79936 4520 79940
rect 34936 79996 35000 80000
rect 34936 79940 34940 79996
rect 34940 79940 34996 79996
rect 34996 79940 35000 79996
rect 34936 79936 35000 79940
rect 35016 79996 35080 80000
rect 35016 79940 35020 79996
rect 35020 79940 35076 79996
rect 35076 79940 35080 79996
rect 35016 79936 35080 79940
rect 35096 79996 35160 80000
rect 35096 79940 35100 79996
rect 35100 79940 35156 79996
rect 35156 79940 35160 79996
rect 35096 79936 35160 79940
rect 35176 79996 35240 80000
rect 35176 79940 35180 79996
rect 35180 79940 35236 79996
rect 35236 79940 35240 79996
rect 35176 79936 35240 79940
rect 65656 79996 65720 80000
rect 65656 79940 65660 79996
rect 65660 79940 65716 79996
rect 65716 79940 65720 79996
rect 65656 79936 65720 79940
rect 65736 79996 65800 80000
rect 65736 79940 65740 79996
rect 65740 79940 65796 79996
rect 65796 79940 65800 79996
rect 65736 79936 65800 79940
rect 65816 79996 65880 80000
rect 65816 79940 65820 79996
rect 65820 79940 65876 79996
rect 65876 79940 65880 79996
rect 65816 79936 65880 79940
rect 65896 79996 65960 80000
rect 65896 79940 65900 79996
rect 65900 79940 65956 79996
rect 65956 79940 65960 79996
rect 65896 79936 65960 79940
rect 96376 79996 96440 80000
rect 96376 79940 96380 79996
rect 96380 79940 96436 79996
rect 96436 79940 96440 79996
rect 96376 79936 96440 79940
rect 96456 79996 96520 80000
rect 96456 79940 96460 79996
rect 96460 79940 96516 79996
rect 96516 79940 96520 79996
rect 96456 79936 96520 79940
rect 96536 79996 96600 80000
rect 96536 79940 96540 79996
rect 96540 79940 96596 79996
rect 96596 79940 96600 79996
rect 96536 79936 96600 79940
rect 96616 79996 96680 80000
rect 96616 79940 96620 79996
rect 96620 79940 96676 79996
rect 96676 79940 96680 79996
rect 96616 79936 96680 79940
rect 4876 79452 4940 79456
rect 4876 79396 4880 79452
rect 4880 79396 4936 79452
rect 4936 79396 4940 79452
rect 4876 79392 4940 79396
rect 4956 79452 5020 79456
rect 4956 79396 4960 79452
rect 4960 79396 5016 79452
rect 5016 79396 5020 79452
rect 4956 79392 5020 79396
rect 5036 79452 5100 79456
rect 5036 79396 5040 79452
rect 5040 79396 5096 79452
rect 5096 79396 5100 79452
rect 5036 79392 5100 79396
rect 5116 79452 5180 79456
rect 5116 79396 5120 79452
rect 5120 79396 5176 79452
rect 5176 79396 5180 79452
rect 5116 79392 5180 79396
rect 35596 79452 35660 79456
rect 35596 79396 35600 79452
rect 35600 79396 35656 79452
rect 35656 79396 35660 79452
rect 35596 79392 35660 79396
rect 35676 79452 35740 79456
rect 35676 79396 35680 79452
rect 35680 79396 35736 79452
rect 35736 79396 35740 79452
rect 35676 79392 35740 79396
rect 35756 79452 35820 79456
rect 35756 79396 35760 79452
rect 35760 79396 35816 79452
rect 35816 79396 35820 79452
rect 35756 79392 35820 79396
rect 35836 79452 35900 79456
rect 35836 79396 35840 79452
rect 35840 79396 35896 79452
rect 35896 79396 35900 79452
rect 35836 79392 35900 79396
rect 66316 79452 66380 79456
rect 66316 79396 66320 79452
rect 66320 79396 66376 79452
rect 66376 79396 66380 79452
rect 66316 79392 66380 79396
rect 66396 79452 66460 79456
rect 66396 79396 66400 79452
rect 66400 79396 66456 79452
rect 66456 79396 66460 79452
rect 66396 79392 66460 79396
rect 66476 79452 66540 79456
rect 66476 79396 66480 79452
rect 66480 79396 66536 79452
rect 66536 79396 66540 79452
rect 66476 79392 66540 79396
rect 66556 79452 66620 79456
rect 66556 79396 66560 79452
rect 66560 79396 66616 79452
rect 66616 79396 66620 79452
rect 66556 79392 66620 79396
rect 97036 79452 97100 79456
rect 97036 79396 97040 79452
rect 97040 79396 97096 79452
rect 97096 79396 97100 79452
rect 97036 79392 97100 79396
rect 97116 79452 97180 79456
rect 97116 79396 97120 79452
rect 97120 79396 97176 79452
rect 97176 79396 97180 79452
rect 97116 79392 97180 79396
rect 97196 79452 97260 79456
rect 97196 79396 97200 79452
rect 97200 79396 97256 79452
rect 97256 79396 97260 79452
rect 97196 79392 97260 79396
rect 97276 79452 97340 79456
rect 97276 79396 97280 79452
rect 97280 79396 97336 79452
rect 97336 79396 97340 79452
rect 97276 79392 97340 79396
rect 4216 78908 4280 78912
rect 4216 78852 4220 78908
rect 4220 78852 4276 78908
rect 4276 78852 4280 78908
rect 4216 78848 4280 78852
rect 4296 78908 4360 78912
rect 4296 78852 4300 78908
rect 4300 78852 4356 78908
rect 4356 78852 4360 78908
rect 4296 78848 4360 78852
rect 4376 78908 4440 78912
rect 4376 78852 4380 78908
rect 4380 78852 4436 78908
rect 4436 78852 4440 78908
rect 4376 78848 4440 78852
rect 4456 78908 4520 78912
rect 4456 78852 4460 78908
rect 4460 78852 4516 78908
rect 4516 78852 4520 78908
rect 4456 78848 4520 78852
rect 34936 78908 35000 78912
rect 34936 78852 34940 78908
rect 34940 78852 34996 78908
rect 34996 78852 35000 78908
rect 34936 78848 35000 78852
rect 35016 78908 35080 78912
rect 35016 78852 35020 78908
rect 35020 78852 35076 78908
rect 35076 78852 35080 78908
rect 35016 78848 35080 78852
rect 35096 78908 35160 78912
rect 35096 78852 35100 78908
rect 35100 78852 35156 78908
rect 35156 78852 35160 78908
rect 35096 78848 35160 78852
rect 35176 78908 35240 78912
rect 35176 78852 35180 78908
rect 35180 78852 35236 78908
rect 35236 78852 35240 78908
rect 35176 78848 35240 78852
rect 65656 78908 65720 78912
rect 65656 78852 65660 78908
rect 65660 78852 65716 78908
rect 65716 78852 65720 78908
rect 65656 78848 65720 78852
rect 65736 78908 65800 78912
rect 65736 78852 65740 78908
rect 65740 78852 65796 78908
rect 65796 78852 65800 78908
rect 65736 78848 65800 78852
rect 65816 78908 65880 78912
rect 65816 78852 65820 78908
rect 65820 78852 65876 78908
rect 65876 78852 65880 78908
rect 65816 78848 65880 78852
rect 65896 78908 65960 78912
rect 65896 78852 65900 78908
rect 65900 78852 65956 78908
rect 65956 78852 65960 78908
rect 65896 78848 65960 78852
rect 96376 78908 96440 78912
rect 96376 78852 96380 78908
rect 96380 78852 96436 78908
rect 96436 78852 96440 78908
rect 96376 78848 96440 78852
rect 96456 78908 96520 78912
rect 96456 78852 96460 78908
rect 96460 78852 96516 78908
rect 96516 78852 96520 78908
rect 96456 78848 96520 78852
rect 96536 78908 96600 78912
rect 96536 78852 96540 78908
rect 96540 78852 96596 78908
rect 96596 78852 96600 78908
rect 96536 78848 96600 78852
rect 96616 78908 96680 78912
rect 96616 78852 96620 78908
rect 96620 78852 96676 78908
rect 96676 78852 96680 78908
rect 96616 78848 96680 78852
rect 4876 78364 4940 78368
rect 4876 78308 4880 78364
rect 4880 78308 4936 78364
rect 4936 78308 4940 78364
rect 4876 78304 4940 78308
rect 4956 78364 5020 78368
rect 4956 78308 4960 78364
rect 4960 78308 5016 78364
rect 5016 78308 5020 78364
rect 4956 78304 5020 78308
rect 5036 78364 5100 78368
rect 5036 78308 5040 78364
rect 5040 78308 5096 78364
rect 5096 78308 5100 78364
rect 5036 78304 5100 78308
rect 5116 78364 5180 78368
rect 5116 78308 5120 78364
rect 5120 78308 5176 78364
rect 5176 78308 5180 78364
rect 5116 78304 5180 78308
rect 35596 78364 35660 78368
rect 35596 78308 35600 78364
rect 35600 78308 35656 78364
rect 35656 78308 35660 78364
rect 35596 78304 35660 78308
rect 35676 78364 35740 78368
rect 35676 78308 35680 78364
rect 35680 78308 35736 78364
rect 35736 78308 35740 78364
rect 35676 78304 35740 78308
rect 35756 78364 35820 78368
rect 35756 78308 35760 78364
rect 35760 78308 35816 78364
rect 35816 78308 35820 78364
rect 35756 78304 35820 78308
rect 35836 78364 35900 78368
rect 35836 78308 35840 78364
rect 35840 78308 35896 78364
rect 35896 78308 35900 78364
rect 35836 78304 35900 78308
rect 66316 78364 66380 78368
rect 66316 78308 66320 78364
rect 66320 78308 66376 78364
rect 66376 78308 66380 78364
rect 66316 78304 66380 78308
rect 66396 78364 66460 78368
rect 66396 78308 66400 78364
rect 66400 78308 66456 78364
rect 66456 78308 66460 78364
rect 66396 78304 66460 78308
rect 66476 78364 66540 78368
rect 66476 78308 66480 78364
rect 66480 78308 66536 78364
rect 66536 78308 66540 78364
rect 66476 78304 66540 78308
rect 66556 78364 66620 78368
rect 66556 78308 66560 78364
rect 66560 78308 66616 78364
rect 66616 78308 66620 78364
rect 66556 78304 66620 78308
rect 97036 78364 97100 78368
rect 97036 78308 97040 78364
rect 97040 78308 97096 78364
rect 97096 78308 97100 78364
rect 97036 78304 97100 78308
rect 97116 78364 97180 78368
rect 97116 78308 97120 78364
rect 97120 78308 97176 78364
rect 97176 78308 97180 78364
rect 97116 78304 97180 78308
rect 97196 78364 97260 78368
rect 97196 78308 97200 78364
rect 97200 78308 97256 78364
rect 97256 78308 97260 78364
rect 97196 78304 97260 78308
rect 97276 78364 97340 78368
rect 97276 78308 97280 78364
rect 97280 78308 97336 78364
rect 97336 78308 97340 78364
rect 97276 78304 97340 78308
rect 4216 77820 4280 77824
rect 4216 77764 4220 77820
rect 4220 77764 4276 77820
rect 4276 77764 4280 77820
rect 4216 77760 4280 77764
rect 4296 77820 4360 77824
rect 4296 77764 4300 77820
rect 4300 77764 4356 77820
rect 4356 77764 4360 77820
rect 4296 77760 4360 77764
rect 4376 77820 4440 77824
rect 4376 77764 4380 77820
rect 4380 77764 4436 77820
rect 4436 77764 4440 77820
rect 4376 77760 4440 77764
rect 4456 77820 4520 77824
rect 4456 77764 4460 77820
rect 4460 77764 4516 77820
rect 4516 77764 4520 77820
rect 4456 77760 4520 77764
rect 34936 77820 35000 77824
rect 34936 77764 34940 77820
rect 34940 77764 34996 77820
rect 34996 77764 35000 77820
rect 34936 77760 35000 77764
rect 35016 77820 35080 77824
rect 35016 77764 35020 77820
rect 35020 77764 35076 77820
rect 35076 77764 35080 77820
rect 35016 77760 35080 77764
rect 35096 77820 35160 77824
rect 35096 77764 35100 77820
rect 35100 77764 35156 77820
rect 35156 77764 35160 77820
rect 35096 77760 35160 77764
rect 35176 77820 35240 77824
rect 35176 77764 35180 77820
rect 35180 77764 35236 77820
rect 35236 77764 35240 77820
rect 35176 77760 35240 77764
rect 65656 77820 65720 77824
rect 65656 77764 65660 77820
rect 65660 77764 65716 77820
rect 65716 77764 65720 77820
rect 65656 77760 65720 77764
rect 65736 77820 65800 77824
rect 65736 77764 65740 77820
rect 65740 77764 65796 77820
rect 65796 77764 65800 77820
rect 65736 77760 65800 77764
rect 65816 77820 65880 77824
rect 65816 77764 65820 77820
rect 65820 77764 65876 77820
rect 65876 77764 65880 77820
rect 65816 77760 65880 77764
rect 65896 77820 65960 77824
rect 65896 77764 65900 77820
rect 65900 77764 65956 77820
rect 65956 77764 65960 77820
rect 65896 77760 65960 77764
rect 96376 77820 96440 77824
rect 96376 77764 96380 77820
rect 96380 77764 96436 77820
rect 96436 77764 96440 77820
rect 96376 77760 96440 77764
rect 96456 77820 96520 77824
rect 96456 77764 96460 77820
rect 96460 77764 96516 77820
rect 96516 77764 96520 77820
rect 96456 77760 96520 77764
rect 96536 77820 96600 77824
rect 96536 77764 96540 77820
rect 96540 77764 96596 77820
rect 96596 77764 96600 77820
rect 96536 77760 96600 77764
rect 96616 77820 96680 77824
rect 96616 77764 96620 77820
rect 96620 77764 96676 77820
rect 96676 77764 96680 77820
rect 96616 77760 96680 77764
rect 4876 77276 4940 77280
rect 4876 77220 4880 77276
rect 4880 77220 4936 77276
rect 4936 77220 4940 77276
rect 4876 77216 4940 77220
rect 4956 77276 5020 77280
rect 4956 77220 4960 77276
rect 4960 77220 5016 77276
rect 5016 77220 5020 77276
rect 4956 77216 5020 77220
rect 5036 77276 5100 77280
rect 5036 77220 5040 77276
rect 5040 77220 5096 77276
rect 5096 77220 5100 77276
rect 5036 77216 5100 77220
rect 5116 77276 5180 77280
rect 5116 77220 5120 77276
rect 5120 77220 5176 77276
rect 5176 77220 5180 77276
rect 5116 77216 5180 77220
rect 35596 77276 35660 77280
rect 35596 77220 35600 77276
rect 35600 77220 35656 77276
rect 35656 77220 35660 77276
rect 35596 77216 35660 77220
rect 35676 77276 35740 77280
rect 35676 77220 35680 77276
rect 35680 77220 35736 77276
rect 35736 77220 35740 77276
rect 35676 77216 35740 77220
rect 35756 77276 35820 77280
rect 35756 77220 35760 77276
rect 35760 77220 35816 77276
rect 35816 77220 35820 77276
rect 35756 77216 35820 77220
rect 35836 77276 35900 77280
rect 35836 77220 35840 77276
rect 35840 77220 35896 77276
rect 35896 77220 35900 77276
rect 35836 77216 35900 77220
rect 66316 77276 66380 77280
rect 66316 77220 66320 77276
rect 66320 77220 66376 77276
rect 66376 77220 66380 77276
rect 66316 77216 66380 77220
rect 66396 77276 66460 77280
rect 66396 77220 66400 77276
rect 66400 77220 66456 77276
rect 66456 77220 66460 77276
rect 66396 77216 66460 77220
rect 66476 77276 66540 77280
rect 66476 77220 66480 77276
rect 66480 77220 66536 77276
rect 66536 77220 66540 77276
rect 66476 77216 66540 77220
rect 66556 77276 66620 77280
rect 66556 77220 66560 77276
rect 66560 77220 66616 77276
rect 66616 77220 66620 77276
rect 66556 77216 66620 77220
rect 97036 77276 97100 77280
rect 97036 77220 97040 77276
rect 97040 77220 97096 77276
rect 97096 77220 97100 77276
rect 97036 77216 97100 77220
rect 97116 77276 97180 77280
rect 97116 77220 97120 77276
rect 97120 77220 97176 77276
rect 97176 77220 97180 77276
rect 97116 77216 97180 77220
rect 97196 77276 97260 77280
rect 97196 77220 97200 77276
rect 97200 77220 97256 77276
rect 97256 77220 97260 77276
rect 97196 77216 97260 77220
rect 97276 77276 97340 77280
rect 97276 77220 97280 77276
rect 97280 77220 97336 77276
rect 97336 77220 97340 77276
rect 97276 77216 97340 77220
rect 45140 77012 45204 77076
rect 4216 76732 4280 76736
rect 4216 76676 4220 76732
rect 4220 76676 4276 76732
rect 4276 76676 4280 76732
rect 4216 76672 4280 76676
rect 4296 76732 4360 76736
rect 4296 76676 4300 76732
rect 4300 76676 4356 76732
rect 4356 76676 4360 76732
rect 4296 76672 4360 76676
rect 4376 76732 4440 76736
rect 4376 76676 4380 76732
rect 4380 76676 4436 76732
rect 4436 76676 4440 76732
rect 4376 76672 4440 76676
rect 4456 76732 4520 76736
rect 4456 76676 4460 76732
rect 4460 76676 4516 76732
rect 4516 76676 4520 76732
rect 4456 76672 4520 76676
rect 34936 76732 35000 76736
rect 34936 76676 34940 76732
rect 34940 76676 34996 76732
rect 34996 76676 35000 76732
rect 34936 76672 35000 76676
rect 35016 76732 35080 76736
rect 35016 76676 35020 76732
rect 35020 76676 35076 76732
rect 35076 76676 35080 76732
rect 35016 76672 35080 76676
rect 35096 76732 35160 76736
rect 35096 76676 35100 76732
rect 35100 76676 35156 76732
rect 35156 76676 35160 76732
rect 35096 76672 35160 76676
rect 35176 76732 35240 76736
rect 35176 76676 35180 76732
rect 35180 76676 35236 76732
rect 35236 76676 35240 76732
rect 35176 76672 35240 76676
rect 65656 76732 65720 76736
rect 65656 76676 65660 76732
rect 65660 76676 65716 76732
rect 65716 76676 65720 76732
rect 65656 76672 65720 76676
rect 65736 76732 65800 76736
rect 65736 76676 65740 76732
rect 65740 76676 65796 76732
rect 65796 76676 65800 76732
rect 65736 76672 65800 76676
rect 65816 76732 65880 76736
rect 65816 76676 65820 76732
rect 65820 76676 65876 76732
rect 65876 76676 65880 76732
rect 65816 76672 65880 76676
rect 65896 76732 65960 76736
rect 65896 76676 65900 76732
rect 65900 76676 65956 76732
rect 65956 76676 65960 76732
rect 65896 76672 65960 76676
rect 96376 76732 96440 76736
rect 96376 76676 96380 76732
rect 96380 76676 96436 76732
rect 96436 76676 96440 76732
rect 96376 76672 96440 76676
rect 96456 76732 96520 76736
rect 96456 76676 96460 76732
rect 96460 76676 96516 76732
rect 96516 76676 96520 76732
rect 96456 76672 96520 76676
rect 96536 76732 96600 76736
rect 96536 76676 96540 76732
rect 96540 76676 96596 76732
rect 96596 76676 96600 76732
rect 96536 76672 96600 76676
rect 96616 76732 96680 76736
rect 96616 76676 96620 76732
rect 96620 76676 96676 76732
rect 96676 76676 96680 76732
rect 96616 76672 96680 76676
rect 37596 76196 37660 76260
rect 4876 76188 4940 76192
rect 4876 76132 4880 76188
rect 4880 76132 4936 76188
rect 4936 76132 4940 76188
rect 4876 76128 4940 76132
rect 4956 76188 5020 76192
rect 4956 76132 4960 76188
rect 4960 76132 5016 76188
rect 5016 76132 5020 76188
rect 4956 76128 5020 76132
rect 5036 76188 5100 76192
rect 5036 76132 5040 76188
rect 5040 76132 5096 76188
rect 5096 76132 5100 76188
rect 5036 76128 5100 76132
rect 5116 76188 5180 76192
rect 5116 76132 5120 76188
rect 5120 76132 5176 76188
rect 5176 76132 5180 76188
rect 5116 76128 5180 76132
rect 35596 76188 35660 76192
rect 35596 76132 35600 76188
rect 35600 76132 35656 76188
rect 35656 76132 35660 76188
rect 35596 76128 35660 76132
rect 35676 76188 35740 76192
rect 35676 76132 35680 76188
rect 35680 76132 35736 76188
rect 35736 76132 35740 76188
rect 35676 76128 35740 76132
rect 35756 76188 35820 76192
rect 35756 76132 35760 76188
rect 35760 76132 35816 76188
rect 35816 76132 35820 76188
rect 35756 76128 35820 76132
rect 35836 76188 35900 76192
rect 35836 76132 35840 76188
rect 35840 76132 35896 76188
rect 35896 76132 35900 76188
rect 35836 76128 35900 76132
rect 66316 76188 66380 76192
rect 66316 76132 66320 76188
rect 66320 76132 66376 76188
rect 66376 76132 66380 76188
rect 66316 76128 66380 76132
rect 66396 76188 66460 76192
rect 66396 76132 66400 76188
rect 66400 76132 66456 76188
rect 66456 76132 66460 76188
rect 66396 76128 66460 76132
rect 66476 76188 66540 76192
rect 66476 76132 66480 76188
rect 66480 76132 66536 76188
rect 66536 76132 66540 76188
rect 66476 76128 66540 76132
rect 66556 76188 66620 76192
rect 66556 76132 66560 76188
rect 66560 76132 66616 76188
rect 66616 76132 66620 76188
rect 66556 76128 66620 76132
rect 97036 76188 97100 76192
rect 97036 76132 97040 76188
rect 97040 76132 97096 76188
rect 97096 76132 97100 76188
rect 97036 76128 97100 76132
rect 97116 76188 97180 76192
rect 97116 76132 97120 76188
rect 97120 76132 97176 76188
rect 97176 76132 97180 76188
rect 97116 76128 97180 76132
rect 97196 76188 97260 76192
rect 97196 76132 97200 76188
rect 97200 76132 97256 76188
rect 97256 76132 97260 76188
rect 97196 76128 97260 76132
rect 97276 76188 97340 76192
rect 97276 76132 97280 76188
rect 97280 76132 97336 76188
rect 97336 76132 97340 76188
rect 97276 76128 97340 76132
rect 42564 75924 42628 75988
rect 50108 75788 50172 75852
rect 4216 75644 4280 75648
rect 4216 75588 4220 75644
rect 4220 75588 4276 75644
rect 4276 75588 4280 75644
rect 4216 75584 4280 75588
rect 4296 75644 4360 75648
rect 4296 75588 4300 75644
rect 4300 75588 4356 75644
rect 4356 75588 4360 75644
rect 4296 75584 4360 75588
rect 4376 75644 4440 75648
rect 4376 75588 4380 75644
rect 4380 75588 4436 75644
rect 4436 75588 4440 75644
rect 4376 75584 4440 75588
rect 4456 75644 4520 75648
rect 4456 75588 4460 75644
rect 4460 75588 4516 75644
rect 4516 75588 4520 75644
rect 4456 75584 4520 75588
rect 34936 75644 35000 75648
rect 34936 75588 34940 75644
rect 34940 75588 34996 75644
rect 34996 75588 35000 75644
rect 34936 75584 35000 75588
rect 35016 75644 35080 75648
rect 35016 75588 35020 75644
rect 35020 75588 35076 75644
rect 35076 75588 35080 75644
rect 35016 75584 35080 75588
rect 35096 75644 35160 75648
rect 35096 75588 35100 75644
rect 35100 75588 35156 75644
rect 35156 75588 35160 75644
rect 35096 75584 35160 75588
rect 35176 75644 35240 75648
rect 35176 75588 35180 75644
rect 35180 75588 35236 75644
rect 35236 75588 35240 75644
rect 35176 75584 35240 75588
rect 65656 75644 65720 75648
rect 65656 75588 65660 75644
rect 65660 75588 65716 75644
rect 65716 75588 65720 75644
rect 65656 75584 65720 75588
rect 65736 75644 65800 75648
rect 65736 75588 65740 75644
rect 65740 75588 65796 75644
rect 65796 75588 65800 75644
rect 65736 75584 65800 75588
rect 65816 75644 65880 75648
rect 65816 75588 65820 75644
rect 65820 75588 65876 75644
rect 65876 75588 65880 75644
rect 65816 75584 65880 75588
rect 65896 75644 65960 75648
rect 65896 75588 65900 75644
rect 65900 75588 65956 75644
rect 65956 75588 65960 75644
rect 65896 75584 65960 75588
rect 96376 75644 96440 75648
rect 96376 75588 96380 75644
rect 96380 75588 96436 75644
rect 96436 75588 96440 75644
rect 96376 75584 96440 75588
rect 96456 75644 96520 75648
rect 96456 75588 96460 75644
rect 96460 75588 96516 75644
rect 96516 75588 96520 75644
rect 96456 75584 96520 75588
rect 96536 75644 96600 75648
rect 96536 75588 96540 75644
rect 96540 75588 96596 75644
rect 96596 75588 96600 75644
rect 96536 75584 96600 75588
rect 96616 75644 96680 75648
rect 96616 75588 96620 75644
rect 96620 75588 96676 75644
rect 96676 75588 96680 75644
rect 96616 75584 96680 75588
rect 4876 75100 4940 75104
rect 4876 75044 4880 75100
rect 4880 75044 4936 75100
rect 4936 75044 4940 75100
rect 4876 75040 4940 75044
rect 4956 75100 5020 75104
rect 4956 75044 4960 75100
rect 4960 75044 5016 75100
rect 5016 75044 5020 75100
rect 4956 75040 5020 75044
rect 5036 75100 5100 75104
rect 5036 75044 5040 75100
rect 5040 75044 5096 75100
rect 5096 75044 5100 75100
rect 5036 75040 5100 75044
rect 5116 75100 5180 75104
rect 5116 75044 5120 75100
rect 5120 75044 5176 75100
rect 5176 75044 5180 75100
rect 5116 75040 5180 75044
rect 35596 75100 35660 75104
rect 35596 75044 35600 75100
rect 35600 75044 35656 75100
rect 35656 75044 35660 75100
rect 35596 75040 35660 75044
rect 35676 75100 35740 75104
rect 35676 75044 35680 75100
rect 35680 75044 35736 75100
rect 35736 75044 35740 75100
rect 35676 75040 35740 75044
rect 35756 75100 35820 75104
rect 35756 75044 35760 75100
rect 35760 75044 35816 75100
rect 35816 75044 35820 75100
rect 35756 75040 35820 75044
rect 35836 75100 35900 75104
rect 35836 75044 35840 75100
rect 35840 75044 35896 75100
rect 35896 75044 35900 75100
rect 35836 75040 35900 75044
rect 66316 75100 66380 75104
rect 66316 75044 66320 75100
rect 66320 75044 66376 75100
rect 66376 75044 66380 75100
rect 66316 75040 66380 75044
rect 66396 75100 66460 75104
rect 66396 75044 66400 75100
rect 66400 75044 66456 75100
rect 66456 75044 66460 75100
rect 66396 75040 66460 75044
rect 66476 75100 66540 75104
rect 66476 75044 66480 75100
rect 66480 75044 66536 75100
rect 66536 75044 66540 75100
rect 66476 75040 66540 75044
rect 66556 75100 66620 75104
rect 66556 75044 66560 75100
rect 66560 75044 66616 75100
rect 66616 75044 66620 75100
rect 66556 75040 66620 75044
rect 97036 75100 97100 75104
rect 97036 75044 97040 75100
rect 97040 75044 97096 75100
rect 97096 75044 97100 75100
rect 97036 75040 97100 75044
rect 97116 75100 97180 75104
rect 97116 75044 97120 75100
rect 97120 75044 97176 75100
rect 97176 75044 97180 75100
rect 97116 75040 97180 75044
rect 97196 75100 97260 75104
rect 97196 75044 97200 75100
rect 97200 75044 97256 75100
rect 97256 75044 97260 75100
rect 97196 75040 97260 75044
rect 97276 75100 97340 75104
rect 97276 75044 97280 75100
rect 97280 75044 97336 75100
rect 97336 75044 97340 75100
rect 97276 75040 97340 75044
rect 40172 74564 40236 74628
rect 52500 74564 52564 74628
rect 4216 74556 4280 74560
rect 4216 74500 4220 74556
rect 4220 74500 4276 74556
rect 4276 74500 4280 74556
rect 4216 74496 4280 74500
rect 4296 74556 4360 74560
rect 4296 74500 4300 74556
rect 4300 74500 4356 74556
rect 4356 74500 4360 74556
rect 4296 74496 4360 74500
rect 4376 74556 4440 74560
rect 4376 74500 4380 74556
rect 4380 74500 4436 74556
rect 4436 74500 4440 74556
rect 4376 74496 4440 74500
rect 4456 74556 4520 74560
rect 4456 74500 4460 74556
rect 4460 74500 4516 74556
rect 4516 74500 4520 74556
rect 4456 74496 4520 74500
rect 34936 74556 35000 74560
rect 34936 74500 34940 74556
rect 34940 74500 34996 74556
rect 34996 74500 35000 74556
rect 34936 74496 35000 74500
rect 35016 74556 35080 74560
rect 35016 74500 35020 74556
rect 35020 74500 35076 74556
rect 35076 74500 35080 74556
rect 35016 74496 35080 74500
rect 35096 74556 35160 74560
rect 35096 74500 35100 74556
rect 35100 74500 35156 74556
rect 35156 74500 35160 74556
rect 35096 74496 35160 74500
rect 35176 74556 35240 74560
rect 35176 74500 35180 74556
rect 35180 74500 35236 74556
rect 35236 74500 35240 74556
rect 35176 74496 35240 74500
rect 65656 74556 65720 74560
rect 65656 74500 65660 74556
rect 65660 74500 65716 74556
rect 65716 74500 65720 74556
rect 65656 74496 65720 74500
rect 65736 74556 65800 74560
rect 65736 74500 65740 74556
rect 65740 74500 65796 74556
rect 65796 74500 65800 74556
rect 65736 74496 65800 74500
rect 65816 74556 65880 74560
rect 65816 74500 65820 74556
rect 65820 74500 65876 74556
rect 65876 74500 65880 74556
rect 65816 74496 65880 74500
rect 65896 74556 65960 74560
rect 65896 74500 65900 74556
rect 65900 74500 65956 74556
rect 65956 74500 65960 74556
rect 65896 74496 65960 74500
rect 96376 74556 96440 74560
rect 96376 74500 96380 74556
rect 96380 74500 96436 74556
rect 96436 74500 96440 74556
rect 96376 74496 96440 74500
rect 96456 74556 96520 74560
rect 96456 74500 96460 74556
rect 96460 74500 96516 74556
rect 96516 74500 96520 74556
rect 96456 74496 96520 74500
rect 96536 74556 96600 74560
rect 96536 74500 96540 74556
rect 96540 74500 96596 74556
rect 96596 74500 96600 74556
rect 96536 74496 96600 74500
rect 96616 74556 96680 74560
rect 96616 74500 96620 74556
rect 96620 74500 96676 74556
rect 96676 74500 96680 74556
rect 96616 74496 96680 74500
rect 4876 74012 4940 74016
rect 4876 73956 4880 74012
rect 4880 73956 4936 74012
rect 4936 73956 4940 74012
rect 4876 73952 4940 73956
rect 4956 74012 5020 74016
rect 4956 73956 4960 74012
rect 4960 73956 5016 74012
rect 5016 73956 5020 74012
rect 4956 73952 5020 73956
rect 5036 74012 5100 74016
rect 5036 73956 5040 74012
rect 5040 73956 5096 74012
rect 5096 73956 5100 74012
rect 5036 73952 5100 73956
rect 5116 74012 5180 74016
rect 5116 73956 5120 74012
rect 5120 73956 5176 74012
rect 5176 73956 5180 74012
rect 5116 73952 5180 73956
rect 35596 74012 35660 74016
rect 35596 73956 35600 74012
rect 35600 73956 35656 74012
rect 35656 73956 35660 74012
rect 35596 73952 35660 73956
rect 35676 74012 35740 74016
rect 35676 73956 35680 74012
rect 35680 73956 35736 74012
rect 35736 73956 35740 74012
rect 35676 73952 35740 73956
rect 35756 74012 35820 74016
rect 35756 73956 35760 74012
rect 35760 73956 35816 74012
rect 35816 73956 35820 74012
rect 35756 73952 35820 73956
rect 35836 74012 35900 74016
rect 35836 73956 35840 74012
rect 35840 73956 35896 74012
rect 35896 73956 35900 74012
rect 35836 73952 35900 73956
rect 66316 74012 66380 74016
rect 66316 73956 66320 74012
rect 66320 73956 66376 74012
rect 66376 73956 66380 74012
rect 66316 73952 66380 73956
rect 66396 74012 66460 74016
rect 66396 73956 66400 74012
rect 66400 73956 66456 74012
rect 66456 73956 66460 74012
rect 66396 73952 66460 73956
rect 66476 74012 66540 74016
rect 66476 73956 66480 74012
rect 66480 73956 66536 74012
rect 66536 73956 66540 74012
rect 66476 73952 66540 73956
rect 66556 74012 66620 74016
rect 66556 73956 66560 74012
rect 66560 73956 66616 74012
rect 66616 73956 66620 74012
rect 66556 73952 66620 73956
rect 97036 74012 97100 74016
rect 97036 73956 97040 74012
rect 97040 73956 97096 74012
rect 97096 73956 97100 74012
rect 97036 73952 97100 73956
rect 97116 74012 97180 74016
rect 97116 73956 97120 74012
rect 97120 73956 97176 74012
rect 97176 73956 97180 74012
rect 97116 73952 97180 73956
rect 97196 74012 97260 74016
rect 97196 73956 97200 74012
rect 97200 73956 97256 74012
rect 97256 73956 97260 74012
rect 97196 73952 97260 73956
rect 97276 74012 97340 74016
rect 97276 73956 97280 74012
rect 97280 73956 97336 74012
rect 97336 73956 97340 74012
rect 97276 73952 97340 73956
rect 55076 73884 55140 73948
rect 4216 73468 4280 73472
rect 4216 73412 4220 73468
rect 4220 73412 4276 73468
rect 4276 73412 4280 73468
rect 4216 73408 4280 73412
rect 4296 73468 4360 73472
rect 4296 73412 4300 73468
rect 4300 73412 4356 73468
rect 4356 73412 4360 73468
rect 4296 73408 4360 73412
rect 4376 73468 4440 73472
rect 4376 73412 4380 73468
rect 4380 73412 4436 73468
rect 4436 73412 4440 73468
rect 4376 73408 4440 73412
rect 4456 73468 4520 73472
rect 4456 73412 4460 73468
rect 4460 73412 4516 73468
rect 4516 73412 4520 73468
rect 4456 73408 4520 73412
rect 34936 73468 35000 73472
rect 34936 73412 34940 73468
rect 34940 73412 34996 73468
rect 34996 73412 35000 73468
rect 34936 73408 35000 73412
rect 35016 73468 35080 73472
rect 35016 73412 35020 73468
rect 35020 73412 35076 73468
rect 35076 73412 35080 73468
rect 35016 73408 35080 73412
rect 35096 73468 35160 73472
rect 35096 73412 35100 73468
rect 35100 73412 35156 73468
rect 35156 73412 35160 73468
rect 35096 73408 35160 73412
rect 35176 73468 35240 73472
rect 35176 73412 35180 73468
rect 35180 73412 35236 73468
rect 35236 73412 35240 73468
rect 35176 73408 35240 73412
rect 65656 73468 65720 73472
rect 65656 73412 65660 73468
rect 65660 73412 65716 73468
rect 65716 73412 65720 73468
rect 65656 73408 65720 73412
rect 65736 73468 65800 73472
rect 65736 73412 65740 73468
rect 65740 73412 65796 73468
rect 65796 73412 65800 73468
rect 65736 73408 65800 73412
rect 65816 73468 65880 73472
rect 65816 73412 65820 73468
rect 65820 73412 65876 73468
rect 65876 73412 65880 73468
rect 65816 73408 65880 73412
rect 65896 73468 65960 73472
rect 65896 73412 65900 73468
rect 65900 73412 65956 73468
rect 65956 73412 65960 73468
rect 65896 73408 65960 73412
rect 96376 73468 96440 73472
rect 96376 73412 96380 73468
rect 96380 73412 96436 73468
rect 96436 73412 96440 73468
rect 96376 73408 96440 73412
rect 96456 73468 96520 73472
rect 96456 73412 96460 73468
rect 96460 73412 96516 73468
rect 96516 73412 96520 73468
rect 96456 73408 96520 73412
rect 96536 73468 96600 73472
rect 96536 73412 96540 73468
rect 96540 73412 96596 73468
rect 96596 73412 96600 73468
rect 96536 73408 96600 73412
rect 96616 73468 96680 73472
rect 96616 73412 96620 73468
rect 96620 73412 96676 73468
rect 96676 73412 96680 73468
rect 96616 73408 96680 73412
rect 4876 72924 4940 72928
rect 4876 72868 4880 72924
rect 4880 72868 4936 72924
rect 4936 72868 4940 72924
rect 4876 72864 4940 72868
rect 4956 72924 5020 72928
rect 4956 72868 4960 72924
rect 4960 72868 5016 72924
rect 5016 72868 5020 72924
rect 4956 72864 5020 72868
rect 5036 72924 5100 72928
rect 5036 72868 5040 72924
rect 5040 72868 5096 72924
rect 5096 72868 5100 72924
rect 5036 72864 5100 72868
rect 5116 72924 5180 72928
rect 5116 72868 5120 72924
rect 5120 72868 5176 72924
rect 5176 72868 5180 72924
rect 5116 72864 5180 72868
rect 35596 72924 35660 72928
rect 35596 72868 35600 72924
rect 35600 72868 35656 72924
rect 35656 72868 35660 72924
rect 35596 72864 35660 72868
rect 35676 72924 35740 72928
rect 35676 72868 35680 72924
rect 35680 72868 35736 72924
rect 35736 72868 35740 72924
rect 35676 72864 35740 72868
rect 35756 72924 35820 72928
rect 35756 72868 35760 72924
rect 35760 72868 35816 72924
rect 35816 72868 35820 72924
rect 35756 72864 35820 72868
rect 35836 72924 35900 72928
rect 35836 72868 35840 72924
rect 35840 72868 35896 72924
rect 35896 72868 35900 72924
rect 35836 72864 35900 72868
rect 66316 72924 66380 72928
rect 66316 72868 66320 72924
rect 66320 72868 66376 72924
rect 66376 72868 66380 72924
rect 66316 72864 66380 72868
rect 66396 72924 66460 72928
rect 66396 72868 66400 72924
rect 66400 72868 66456 72924
rect 66456 72868 66460 72924
rect 66396 72864 66460 72868
rect 66476 72924 66540 72928
rect 66476 72868 66480 72924
rect 66480 72868 66536 72924
rect 66536 72868 66540 72924
rect 66476 72864 66540 72868
rect 66556 72924 66620 72928
rect 66556 72868 66560 72924
rect 66560 72868 66616 72924
rect 66616 72868 66620 72924
rect 66556 72864 66620 72868
rect 97036 72924 97100 72928
rect 97036 72868 97040 72924
rect 97040 72868 97096 72924
rect 97096 72868 97100 72924
rect 97036 72864 97100 72868
rect 97116 72924 97180 72928
rect 97116 72868 97120 72924
rect 97120 72868 97176 72924
rect 97176 72868 97180 72924
rect 97116 72864 97180 72868
rect 97196 72924 97260 72928
rect 97196 72868 97200 72924
rect 97200 72868 97256 72924
rect 97256 72868 97260 72924
rect 97196 72864 97260 72868
rect 97276 72924 97340 72928
rect 97276 72868 97280 72924
rect 97280 72868 97336 72924
rect 97336 72868 97340 72924
rect 97276 72864 97340 72868
rect 4216 72380 4280 72384
rect 4216 72324 4220 72380
rect 4220 72324 4276 72380
rect 4276 72324 4280 72380
rect 4216 72320 4280 72324
rect 4296 72380 4360 72384
rect 4296 72324 4300 72380
rect 4300 72324 4356 72380
rect 4356 72324 4360 72380
rect 4296 72320 4360 72324
rect 4376 72380 4440 72384
rect 4376 72324 4380 72380
rect 4380 72324 4436 72380
rect 4436 72324 4440 72380
rect 4376 72320 4440 72324
rect 4456 72380 4520 72384
rect 4456 72324 4460 72380
rect 4460 72324 4516 72380
rect 4516 72324 4520 72380
rect 4456 72320 4520 72324
rect 34936 72380 35000 72384
rect 34936 72324 34940 72380
rect 34940 72324 34996 72380
rect 34996 72324 35000 72380
rect 34936 72320 35000 72324
rect 35016 72380 35080 72384
rect 35016 72324 35020 72380
rect 35020 72324 35076 72380
rect 35076 72324 35080 72380
rect 35016 72320 35080 72324
rect 35096 72380 35160 72384
rect 35096 72324 35100 72380
rect 35100 72324 35156 72380
rect 35156 72324 35160 72380
rect 35096 72320 35160 72324
rect 35176 72380 35240 72384
rect 35176 72324 35180 72380
rect 35180 72324 35236 72380
rect 35236 72324 35240 72380
rect 35176 72320 35240 72324
rect 65656 72380 65720 72384
rect 65656 72324 65660 72380
rect 65660 72324 65716 72380
rect 65716 72324 65720 72380
rect 65656 72320 65720 72324
rect 65736 72380 65800 72384
rect 65736 72324 65740 72380
rect 65740 72324 65796 72380
rect 65796 72324 65800 72380
rect 65736 72320 65800 72324
rect 65816 72380 65880 72384
rect 65816 72324 65820 72380
rect 65820 72324 65876 72380
rect 65876 72324 65880 72380
rect 65816 72320 65880 72324
rect 65896 72380 65960 72384
rect 65896 72324 65900 72380
rect 65900 72324 65956 72380
rect 65956 72324 65960 72380
rect 65896 72320 65960 72324
rect 96376 72380 96440 72384
rect 96376 72324 96380 72380
rect 96380 72324 96436 72380
rect 96436 72324 96440 72380
rect 96376 72320 96440 72324
rect 96456 72380 96520 72384
rect 96456 72324 96460 72380
rect 96460 72324 96516 72380
rect 96516 72324 96520 72380
rect 96456 72320 96520 72324
rect 96536 72380 96600 72384
rect 96536 72324 96540 72380
rect 96540 72324 96596 72380
rect 96596 72324 96600 72380
rect 96536 72320 96600 72324
rect 96616 72380 96680 72384
rect 96616 72324 96620 72380
rect 96620 72324 96676 72380
rect 96676 72324 96680 72380
rect 96616 72320 96680 72324
rect 47532 71844 47596 71908
rect 4876 71836 4940 71840
rect 4876 71780 4880 71836
rect 4880 71780 4936 71836
rect 4936 71780 4940 71836
rect 4876 71776 4940 71780
rect 4956 71836 5020 71840
rect 4956 71780 4960 71836
rect 4960 71780 5016 71836
rect 5016 71780 5020 71836
rect 4956 71776 5020 71780
rect 5036 71836 5100 71840
rect 5036 71780 5040 71836
rect 5040 71780 5096 71836
rect 5096 71780 5100 71836
rect 5036 71776 5100 71780
rect 5116 71836 5180 71840
rect 5116 71780 5120 71836
rect 5120 71780 5176 71836
rect 5176 71780 5180 71836
rect 5116 71776 5180 71780
rect 35596 71836 35660 71840
rect 35596 71780 35600 71836
rect 35600 71780 35656 71836
rect 35656 71780 35660 71836
rect 35596 71776 35660 71780
rect 35676 71836 35740 71840
rect 35676 71780 35680 71836
rect 35680 71780 35736 71836
rect 35736 71780 35740 71836
rect 35676 71776 35740 71780
rect 35756 71836 35820 71840
rect 35756 71780 35760 71836
rect 35760 71780 35816 71836
rect 35816 71780 35820 71836
rect 35756 71776 35820 71780
rect 35836 71836 35900 71840
rect 35836 71780 35840 71836
rect 35840 71780 35896 71836
rect 35896 71780 35900 71836
rect 35836 71776 35900 71780
rect 66316 71836 66380 71840
rect 66316 71780 66320 71836
rect 66320 71780 66376 71836
rect 66376 71780 66380 71836
rect 66316 71776 66380 71780
rect 66396 71836 66460 71840
rect 66396 71780 66400 71836
rect 66400 71780 66456 71836
rect 66456 71780 66460 71836
rect 66396 71776 66460 71780
rect 66476 71836 66540 71840
rect 66476 71780 66480 71836
rect 66480 71780 66536 71836
rect 66536 71780 66540 71836
rect 66476 71776 66540 71780
rect 66556 71836 66620 71840
rect 66556 71780 66560 71836
rect 66560 71780 66616 71836
rect 66616 71780 66620 71836
rect 66556 71776 66620 71780
rect 97036 71836 97100 71840
rect 97036 71780 97040 71836
rect 97040 71780 97096 71836
rect 97096 71780 97100 71836
rect 97036 71776 97100 71780
rect 97116 71836 97180 71840
rect 97116 71780 97120 71836
rect 97120 71780 97176 71836
rect 97176 71780 97180 71836
rect 97116 71776 97180 71780
rect 97196 71836 97260 71840
rect 97196 71780 97200 71836
rect 97200 71780 97256 71836
rect 97256 71780 97260 71836
rect 97196 71776 97260 71780
rect 97276 71836 97340 71840
rect 97276 71780 97280 71836
rect 97280 71780 97336 71836
rect 97336 71780 97340 71836
rect 97276 71776 97340 71780
rect 4216 71292 4280 71296
rect 4216 71236 4220 71292
rect 4220 71236 4276 71292
rect 4276 71236 4280 71292
rect 4216 71232 4280 71236
rect 4296 71292 4360 71296
rect 4296 71236 4300 71292
rect 4300 71236 4356 71292
rect 4356 71236 4360 71292
rect 4296 71232 4360 71236
rect 4376 71292 4440 71296
rect 4376 71236 4380 71292
rect 4380 71236 4436 71292
rect 4436 71236 4440 71292
rect 4376 71232 4440 71236
rect 4456 71292 4520 71296
rect 4456 71236 4460 71292
rect 4460 71236 4516 71292
rect 4516 71236 4520 71292
rect 4456 71232 4520 71236
rect 34936 71292 35000 71296
rect 34936 71236 34940 71292
rect 34940 71236 34996 71292
rect 34996 71236 35000 71292
rect 34936 71232 35000 71236
rect 35016 71292 35080 71296
rect 35016 71236 35020 71292
rect 35020 71236 35076 71292
rect 35076 71236 35080 71292
rect 35016 71232 35080 71236
rect 35096 71292 35160 71296
rect 35096 71236 35100 71292
rect 35100 71236 35156 71292
rect 35156 71236 35160 71292
rect 35096 71232 35160 71236
rect 35176 71292 35240 71296
rect 35176 71236 35180 71292
rect 35180 71236 35236 71292
rect 35236 71236 35240 71292
rect 35176 71232 35240 71236
rect 65656 71292 65720 71296
rect 65656 71236 65660 71292
rect 65660 71236 65716 71292
rect 65716 71236 65720 71292
rect 65656 71232 65720 71236
rect 65736 71292 65800 71296
rect 65736 71236 65740 71292
rect 65740 71236 65796 71292
rect 65796 71236 65800 71292
rect 65736 71232 65800 71236
rect 65816 71292 65880 71296
rect 65816 71236 65820 71292
rect 65820 71236 65876 71292
rect 65876 71236 65880 71292
rect 65816 71232 65880 71236
rect 65896 71292 65960 71296
rect 65896 71236 65900 71292
rect 65900 71236 65956 71292
rect 65956 71236 65960 71292
rect 65896 71232 65960 71236
rect 96376 71292 96440 71296
rect 96376 71236 96380 71292
rect 96380 71236 96436 71292
rect 96436 71236 96440 71292
rect 96376 71232 96440 71236
rect 96456 71292 96520 71296
rect 96456 71236 96460 71292
rect 96460 71236 96516 71292
rect 96516 71236 96520 71292
rect 96456 71232 96520 71236
rect 96536 71292 96600 71296
rect 96536 71236 96540 71292
rect 96540 71236 96596 71292
rect 96596 71236 96600 71292
rect 96536 71232 96600 71236
rect 96616 71292 96680 71296
rect 96616 71236 96620 71292
rect 96620 71236 96676 71292
rect 96676 71236 96680 71292
rect 96616 71232 96680 71236
rect 4876 70748 4940 70752
rect 4876 70692 4880 70748
rect 4880 70692 4936 70748
rect 4936 70692 4940 70748
rect 4876 70688 4940 70692
rect 4956 70748 5020 70752
rect 4956 70692 4960 70748
rect 4960 70692 5016 70748
rect 5016 70692 5020 70748
rect 4956 70688 5020 70692
rect 5036 70748 5100 70752
rect 5036 70692 5040 70748
rect 5040 70692 5096 70748
rect 5096 70692 5100 70748
rect 5036 70688 5100 70692
rect 5116 70748 5180 70752
rect 5116 70692 5120 70748
rect 5120 70692 5176 70748
rect 5176 70692 5180 70748
rect 5116 70688 5180 70692
rect 35596 70748 35660 70752
rect 35596 70692 35600 70748
rect 35600 70692 35656 70748
rect 35656 70692 35660 70748
rect 35596 70688 35660 70692
rect 35676 70748 35740 70752
rect 35676 70692 35680 70748
rect 35680 70692 35736 70748
rect 35736 70692 35740 70748
rect 35676 70688 35740 70692
rect 35756 70748 35820 70752
rect 35756 70692 35760 70748
rect 35760 70692 35816 70748
rect 35816 70692 35820 70748
rect 35756 70688 35820 70692
rect 35836 70748 35900 70752
rect 35836 70692 35840 70748
rect 35840 70692 35896 70748
rect 35896 70692 35900 70748
rect 35836 70688 35900 70692
rect 66316 70748 66380 70752
rect 66316 70692 66320 70748
rect 66320 70692 66376 70748
rect 66376 70692 66380 70748
rect 66316 70688 66380 70692
rect 66396 70748 66460 70752
rect 66396 70692 66400 70748
rect 66400 70692 66456 70748
rect 66456 70692 66460 70748
rect 66396 70688 66460 70692
rect 66476 70748 66540 70752
rect 66476 70692 66480 70748
rect 66480 70692 66536 70748
rect 66536 70692 66540 70748
rect 66476 70688 66540 70692
rect 66556 70748 66620 70752
rect 66556 70692 66560 70748
rect 66560 70692 66616 70748
rect 66616 70692 66620 70748
rect 66556 70688 66620 70692
rect 97036 70748 97100 70752
rect 97036 70692 97040 70748
rect 97040 70692 97096 70748
rect 97096 70692 97100 70748
rect 97036 70688 97100 70692
rect 97116 70748 97180 70752
rect 97116 70692 97120 70748
rect 97120 70692 97176 70748
rect 97176 70692 97180 70748
rect 97116 70688 97180 70692
rect 97196 70748 97260 70752
rect 97196 70692 97200 70748
rect 97200 70692 97256 70748
rect 97256 70692 97260 70748
rect 97196 70688 97260 70692
rect 97276 70748 97340 70752
rect 97276 70692 97280 70748
rect 97280 70692 97336 70748
rect 97336 70692 97340 70748
rect 97276 70688 97340 70692
rect 4216 70204 4280 70208
rect 4216 70148 4220 70204
rect 4220 70148 4276 70204
rect 4276 70148 4280 70204
rect 4216 70144 4280 70148
rect 4296 70204 4360 70208
rect 4296 70148 4300 70204
rect 4300 70148 4356 70204
rect 4356 70148 4360 70204
rect 4296 70144 4360 70148
rect 4376 70204 4440 70208
rect 4376 70148 4380 70204
rect 4380 70148 4436 70204
rect 4436 70148 4440 70204
rect 4376 70144 4440 70148
rect 4456 70204 4520 70208
rect 4456 70148 4460 70204
rect 4460 70148 4516 70204
rect 4516 70148 4520 70204
rect 4456 70144 4520 70148
rect 34936 70204 35000 70208
rect 34936 70148 34940 70204
rect 34940 70148 34996 70204
rect 34996 70148 35000 70204
rect 34936 70144 35000 70148
rect 35016 70204 35080 70208
rect 35016 70148 35020 70204
rect 35020 70148 35076 70204
rect 35076 70148 35080 70204
rect 35016 70144 35080 70148
rect 35096 70204 35160 70208
rect 35096 70148 35100 70204
rect 35100 70148 35156 70204
rect 35156 70148 35160 70204
rect 35096 70144 35160 70148
rect 35176 70204 35240 70208
rect 35176 70148 35180 70204
rect 35180 70148 35236 70204
rect 35236 70148 35240 70204
rect 35176 70144 35240 70148
rect 65656 70204 65720 70208
rect 65656 70148 65660 70204
rect 65660 70148 65716 70204
rect 65716 70148 65720 70204
rect 65656 70144 65720 70148
rect 65736 70204 65800 70208
rect 65736 70148 65740 70204
rect 65740 70148 65796 70204
rect 65796 70148 65800 70204
rect 65736 70144 65800 70148
rect 65816 70204 65880 70208
rect 65816 70148 65820 70204
rect 65820 70148 65876 70204
rect 65876 70148 65880 70204
rect 65816 70144 65880 70148
rect 65896 70204 65960 70208
rect 65896 70148 65900 70204
rect 65900 70148 65956 70204
rect 65956 70148 65960 70204
rect 65896 70144 65960 70148
rect 96376 70204 96440 70208
rect 96376 70148 96380 70204
rect 96380 70148 96436 70204
rect 96436 70148 96440 70204
rect 96376 70144 96440 70148
rect 96456 70204 96520 70208
rect 96456 70148 96460 70204
rect 96460 70148 96516 70204
rect 96516 70148 96520 70204
rect 96456 70144 96520 70148
rect 96536 70204 96600 70208
rect 96536 70148 96540 70204
rect 96540 70148 96596 70204
rect 96596 70148 96600 70204
rect 96536 70144 96600 70148
rect 96616 70204 96680 70208
rect 96616 70148 96620 70204
rect 96620 70148 96676 70204
rect 96676 70148 96680 70204
rect 96616 70144 96680 70148
rect 4876 69660 4940 69664
rect 4876 69604 4880 69660
rect 4880 69604 4936 69660
rect 4936 69604 4940 69660
rect 4876 69600 4940 69604
rect 4956 69660 5020 69664
rect 4956 69604 4960 69660
rect 4960 69604 5016 69660
rect 5016 69604 5020 69660
rect 4956 69600 5020 69604
rect 5036 69660 5100 69664
rect 5036 69604 5040 69660
rect 5040 69604 5096 69660
rect 5096 69604 5100 69660
rect 5036 69600 5100 69604
rect 5116 69660 5180 69664
rect 5116 69604 5120 69660
rect 5120 69604 5176 69660
rect 5176 69604 5180 69660
rect 5116 69600 5180 69604
rect 35596 69660 35660 69664
rect 35596 69604 35600 69660
rect 35600 69604 35656 69660
rect 35656 69604 35660 69660
rect 35596 69600 35660 69604
rect 35676 69660 35740 69664
rect 35676 69604 35680 69660
rect 35680 69604 35736 69660
rect 35736 69604 35740 69660
rect 35676 69600 35740 69604
rect 35756 69660 35820 69664
rect 35756 69604 35760 69660
rect 35760 69604 35816 69660
rect 35816 69604 35820 69660
rect 35756 69600 35820 69604
rect 35836 69660 35900 69664
rect 35836 69604 35840 69660
rect 35840 69604 35896 69660
rect 35896 69604 35900 69660
rect 35836 69600 35900 69604
rect 66316 69660 66380 69664
rect 66316 69604 66320 69660
rect 66320 69604 66376 69660
rect 66376 69604 66380 69660
rect 66316 69600 66380 69604
rect 66396 69660 66460 69664
rect 66396 69604 66400 69660
rect 66400 69604 66456 69660
rect 66456 69604 66460 69660
rect 66396 69600 66460 69604
rect 66476 69660 66540 69664
rect 66476 69604 66480 69660
rect 66480 69604 66536 69660
rect 66536 69604 66540 69660
rect 66476 69600 66540 69604
rect 66556 69660 66620 69664
rect 66556 69604 66560 69660
rect 66560 69604 66616 69660
rect 66616 69604 66620 69660
rect 66556 69600 66620 69604
rect 97036 69660 97100 69664
rect 97036 69604 97040 69660
rect 97040 69604 97096 69660
rect 97096 69604 97100 69660
rect 97036 69600 97100 69604
rect 97116 69660 97180 69664
rect 97116 69604 97120 69660
rect 97120 69604 97176 69660
rect 97176 69604 97180 69660
rect 97116 69600 97180 69604
rect 97196 69660 97260 69664
rect 97196 69604 97200 69660
rect 97200 69604 97256 69660
rect 97256 69604 97260 69660
rect 97196 69600 97260 69604
rect 97276 69660 97340 69664
rect 97276 69604 97280 69660
rect 97280 69604 97336 69660
rect 97336 69604 97340 69660
rect 97276 69600 97340 69604
rect 4216 69116 4280 69120
rect 4216 69060 4220 69116
rect 4220 69060 4276 69116
rect 4276 69060 4280 69116
rect 4216 69056 4280 69060
rect 4296 69116 4360 69120
rect 4296 69060 4300 69116
rect 4300 69060 4356 69116
rect 4356 69060 4360 69116
rect 4296 69056 4360 69060
rect 4376 69116 4440 69120
rect 4376 69060 4380 69116
rect 4380 69060 4436 69116
rect 4436 69060 4440 69116
rect 4376 69056 4440 69060
rect 4456 69116 4520 69120
rect 4456 69060 4460 69116
rect 4460 69060 4516 69116
rect 4516 69060 4520 69116
rect 4456 69056 4520 69060
rect 34936 69116 35000 69120
rect 34936 69060 34940 69116
rect 34940 69060 34996 69116
rect 34996 69060 35000 69116
rect 34936 69056 35000 69060
rect 35016 69116 35080 69120
rect 35016 69060 35020 69116
rect 35020 69060 35076 69116
rect 35076 69060 35080 69116
rect 35016 69056 35080 69060
rect 35096 69116 35160 69120
rect 35096 69060 35100 69116
rect 35100 69060 35156 69116
rect 35156 69060 35160 69116
rect 35096 69056 35160 69060
rect 35176 69116 35240 69120
rect 35176 69060 35180 69116
rect 35180 69060 35236 69116
rect 35236 69060 35240 69116
rect 35176 69056 35240 69060
rect 65656 69116 65720 69120
rect 65656 69060 65660 69116
rect 65660 69060 65716 69116
rect 65716 69060 65720 69116
rect 65656 69056 65720 69060
rect 65736 69116 65800 69120
rect 65736 69060 65740 69116
rect 65740 69060 65796 69116
rect 65796 69060 65800 69116
rect 65736 69056 65800 69060
rect 65816 69116 65880 69120
rect 65816 69060 65820 69116
rect 65820 69060 65876 69116
rect 65876 69060 65880 69116
rect 65816 69056 65880 69060
rect 65896 69116 65960 69120
rect 65896 69060 65900 69116
rect 65900 69060 65956 69116
rect 65956 69060 65960 69116
rect 65896 69056 65960 69060
rect 96376 69116 96440 69120
rect 96376 69060 96380 69116
rect 96380 69060 96436 69116
rect 96436 69060 96440 69116
rect 96376 69056 96440 69060
rect 96456 69116 96520 69120
rect 96456 69060 96460 69116
rect 96460 69060 96516 69116
rect 96516 69060 96520 69116
rect 96456 69056 96520 69060
rect 96536 69116 96600 69120
rect 96536 69060 96540 69116
rect 96540 69060 96596 69116
rect 96596 69060 96600 69116
rect 96536 69056 96600 69060
rect 96616 69116 96680 69120
rect 96616 69060 96620 69116
rect 96620 69060 96676 69116
rect 96676 69060 96680 69116
rect 96616 69056 96680 69060
rect 4876 68572 4940 68576
rect 4876 68516 4880 68572
rect 4880 68516 4936 68572
rect 4936 68516 4940 68572
rect 4876 68512 4940 68516
rect 4956 68572 5020 68576
rect 4956 68516 4960 68572
rect 4960 68516 5016 68572
rect 5016 68516 5020 68572
rect 4956 68512 5020 68516
rect 5036 68572 5100 68576
rect 5036 68516 5040 68572
rect 5040 68516 5096 68572
rect 5096 68516 5100 68572
rect 5036 68512 5100 68516
rect 5116 68572 5180 68576
rect 5116 68516 5120 68572
rect 5120 68516 5176 68572
rect 5176 68516 5180 68572
rect 5116 68512 5180 68516
rect 35596 68572 35660 68576
rect 35596 68516 35600 68572
rect 35600 68516 35656 68572
rect 35656 68516 35660 68572
rect 35596 68512 35660 68516
rect 35676 68572 35740 68576
rect 35676 68516 35680 68572
rect 35680 68516 35736 68572
rect 35736 68516 35740 68572
rect 35676 68512 35740 68516
rect 35756 68572 35820 68576
rect 35756 68516 35760 68572
rect 35760 68516 35816 68572
rect 35816 68516 35820 68572
rect 35756 68512 35820 68516
rect 35836 68572 35900 68576
rect 35836 68516 35840 68572
rect 35840 68516 35896 68572
rect 35896 68516 35900 68572
rect 35836 68512 35900 68516
rect 66316 68572 66380 68576
rect 66316 68516 66320 68572
rect 66320 68516 66376 68572
rect 66376 68516 66380 68572
rect 66316 68512 66380 68516
rect 66396 68572 66460 68576
rect 66396 68516 66400 68572
rect 66400 68516 66456 68572
rect 66456 68516 66460 68572
rect 66396 68512 66460 68516
rect 66476 68572 66540 68576
rect 66476 68516 66480 68572
rect 66480 68516 66536 68572
rect 66536 68516 66540 68572
rect 66476 68512 66540 68516
rect 66556 68572 66620 68576
rect 66556 68516 66560 68572
rect 66560 68516 66616 68572
rect 66616 68516 66620 68572
rect 66556 68512 66620 68516
rect 97036 68572 97100 68576
rect 97036 68516 97040 68572
rect 97040 68516 97096 68572
rect 97096 68516 97100 68572
rect 97036 68512 97100 68516
rect 97116 68572 97180 68576
rect 97116 68516 97120 68572
rect 97120 68516 97176 68572
rect 97176 68516 97180 68572
rect 97116 68512 97180 68516
rect 97196 68572 97260 68576
rect 97196 68516 97200 68572
rect 97200 68516 97256 68572
rect 97256 68516 97260 68572
rect 97196 68512 97260 68516
rect 97276 68572 97340 68576
rect 97276 68516 97280 68572
rect 97280 68516 97336 68572
rect 97336 68516 97340 68572
rect 97276 68512 97340 68516
rect 4216 68028 4280 68032
rect 4216 67972 4220 68028
rect 4220 67972 4276 68028
rect 4276 67972 4280 68028
rect 4216 67968 4280 67972
rect 4296 68028 4360 68032
rect 4296 67972 4300 68028
rect 4300 67972 4356 68028
rect 4356 67972 4360 68028
rect 4296 67968 4360 67972
rect 4376 68028 4440 68032
rect 4376 67972 4380 68028
rect 4380 67972 4436 68028
rect 4436 67972 4440 68028
rect 4376 67968 4440 67972
rect 4456 68028 4520 68032
rect 4456 67972 4460 68028
rect 4460 67972 4516 68028
rect 4516 67972 4520 68028
rect 4456 67968 4520 67972
rect 34936 68028 35000 68032
rect 34936 67972 34940 68028
rect 34940 67972 34996 68028
rect 34996 67972 35000 68028
rect 34936 67968 35000 67972
rect 35016 68028 35080 68032
rect 35016 67972 35020 68028
rect 35020 67972 35076 68028
rect 35076 67972 35080 68028
rect 35016 67968 35080 67972
rect 35096 68028 35160 68032
rect 35096 67972 35100 68028
rect 35100 67972 35156 68028
rect 35156 67972 35160 68028
rect 35096 67968 35160 67972
rect 35176 68028 35240 68032
rect 35176 67972 35180 68028
rect 35180 67972 35236 68028
rect 35236 67972 35240 68028
rect 35176 67968 35240 67972
rect 65656 68028 65720 68032
rect 65656 67972 65660 68028
rect 65660 67972 65716 68028
rect 65716 67972 65720 68028
rect 65656 67968 65720 67972
rect 65736 68028 65800 68032
rect 65736 67972 65740 68028
rect 65740 67972 65796 68028
rect 65796 67972 65800 68028
rect 65736 67968 65800 67972
rect 65816 68028 65880 68032
rect 65816 67972 65820 68028
rect 65820 67972 65876 68028
rect 65876 67972 65880 68028
rect 65816 67968 65880 67972
rect 65896 68028 65960 68032
rect 65896 67972 65900 68028
rect 65900 67972 65956 68028
rect 65956 67972 65960 68028
rect 65896 67968 65960 67972
rect 96376 68028 96440 68032
rect 96376 67972 96380 68028
rect 96380 67972 96436 68028
rect 96436 67972 96440 68028
rect 96376 67968 96440 67972
rect 96456 68028 96520 68032
rect 96456 67972 96460 68028
rect 96460 67972 96516 68028
rect 96516 67972 96520 68028
rect 96456 67968 96520 67972
rect 96536 68028 96600 68032
rect 96536 67972 96540 68028
rect 96540 67972 96596 68028
rect 96596 67972 96600 68028
rect 96536 67968 96600 67972
rect 96616 68028 96680 68032
rect 96616 67972 96620 68028
rect 96620 67972 96676 68028
rect 96676 67972 96680 68028
rect 96616 67968 96680 67972
rect 4876 67484 4940 67488
rect 4876 67428 4880 67484
rect 4880 67428 4936 67484
rect 4936 67428 4940 67484
rect 4876 67424 4940 67428
rect 4956 67484 5020 67488
rect 4956 67428 4960 67484
rect 4960 67428 5016 67484
rect 5016 67428 5020 67484
rect 4956 67424 5020 67428
rect 5036 67484 5100 67488
rect 5036 67428 5040 67484
rect 5040 67428 5096 67484
rect 5096 67428 5100 67484
rect 5036 67424 5100 67428
rect 5116 67484 5180 67488
rect 5116 67428 5120 67484
rect 5120 67428 5176 67484
rect 5176 67428 5180 67484
rect 5116 67424 5180 67428
rect 35596 67484 35660 67488
rect 35596 67428 35600 67484
rect 35600 67428 35656 67484
rect 35656 67428 35660 67484
rect 35596 67424 35660 67428
rect 35676 67484 35740 67488
rect 35676 67428 35680 67484
rect 35680 67428 35736 67484
rect 35736 67428 35740 67484
rect 35676 67424 35740 67428
rect 35756 67484 35820 67488
rect 35756 67428 35760 67484
rect 35760 67428 35816 67484
rect 35816 67428 35820 67484
rect 35756 67424 35820 67428
rect 35836 67484 35900 67488
rect 35836 67428 35840 67484
rect 35840 67428 35896 67484
rect 35896 67428 35900 67484
rect 35836 67424 35900 67428
rect 66316 67484 66380 67488
rect 66316 67428 66320 67484
rect 66320 67428 66376 67484
rect 66376 67428 66380 67484
rect 66316 67424 66380 67428
rect 66396 67484 66460 67488
rect 66396 67428 66400 67484
rect 66400 67428 66456 67484
rect 66456 67428 66460 67484
rect 66396 67424 66460 67428
rect 66476 67484 66540 67488
rect 66476 67428 66480 67484
rect 66480 67428 66536 67484
rect 66536 67428 66540 67484
rect 66476 67424 66540 67428
rect 66556 67484 66620 67488
rect 66556 67428 66560 67484
rect 66560 67428 66616 67484
rect 66616 67428 66620 67484
rect 66556 67424 66620 67428
rect 97036 67484 97100 67488
rect 97036 67428 97040 67484
rect 97040 67428 97096 67484
rect 97096 67428 97100 67484
rect 97036 67424 97100 67428
rect 97116 67484 97180 67488
rect 97116 67428 97120 67484
rect 97120 67428 97176 67484
rect 97176 67428 97180 67484
rect 97116 67424 97180 67428
rect 97196 67484 97260 67488
rect 97196 67428 97200 67484
rect 97200 67428 97256 67484
rect 97256 67428 97260 67484
rect 97196 67424 97260 67428
rect 97276 67484 97340 67488
rect 97276 67428 97280 67484
rect 97280 67428 97336 67484
rect 97336 67428 97340 67484
rect 97276 67424 97340 67428
rect 4216 66940 4280 66944
rect 4216 66884 4220 66940
rect 4220 66884 4276 66940
rect 4276 66884 4280 66940
rect 4216 66880 4280 66884
rect 4296 66940 4360 66944
rect 4296 66884 4300 66940
rect 4300 66884 4356 66940
rect 4356 66884 4360 66940
rect 4296 66880 4360 66884
rect 4376 66940 4440 66944
rect 4376 66884 4380 66940
rect 4380 66884 4436 66940
rect 4436 66884 4440 66940
rect 4376 66880 4440 66884
rect 4456 66940 4520 66944
rect 4456 66884 4460 66940
rect 4460 66884 4516 66940
rect 4516 66884 4520 66940
rect 4456 66880 4520 66884
rect 34936 66940 35000 66944
rect 34936 66884 34940 66940
rect 34940 66884 34996 66940
rect 34996 66884 35000 66940
rect 34936 66880 35000 66884
rect 35016 66940 35080 66944
rect 35016 66884 35020 66940
rect 35020 66884 35076 66940
rect 35076 66884 35080 66940
rect 35016 66880 35080 66884
rect 35096 66940 35160 66944
rect 35096 66884 35100 66940
rect 35100 66884 35156 66940
rect 35156 66884 35160 66940
rect 35096 66880 35160 66884
rect 35176 66940 35240 66944
rect 35176 66884 35180 66940
rect 35180 66884 35236 66940
rect 35236 66884 35240 66940
rect 35176 66880 35240 66884
rect 65656 66940 65720 66944
rect 65656 66884 65660 66940
rect 65660 66884 65716 66940
rect 65716 66884 65720 66940
rect 65656 66880 65720 66884
rect 65736 66940 65800 66944
rect 65736 66884 65740 66940
rect 65740 66884 65796 66940
rect 65796 66884 65800 66940
rect 65736 66880 65800 66884
rect 65816 66940 65880 66944
rect 65816 66884 65820 66940
rect 65820 66884 65876 66940
rect 65876 66884 65880 66940
rect 65816 66880 65880 66884
rect 65896 66940 65960 66944
rect 65896 66884 65900 66940
rect 65900 66884 65956 66940
rect 65956 66884 65960 66940
rect 65896 66880 65960 66884
rect 96376 66940 96440 66944
rect 96376 66884 96380 66940
rect 96380 66884 96436 66940
rect 96436 66884 96440 66940
rect 96376 66880 96440 66884
rect 96456 66940 96520 66944
rect 96456 66884 96460 66940
rect 96460 66884 96516 66940
rect 96516 66884 96520 66940
rect 96456 66880 96520 66884
rect 96536 66940 96600 66944
rect 96536 66884 96540 66940
rect 96540 66884 96596 66940
rect 96596 66884 96600 66940
rect 96536 66880 96600 66884
rect 96616 66940 96680 66944
rect 96616 66884 96620 66940
rect 96620 66884 96676 66940
rect 96676 66884 96680 66940
rect 96616 66880 96680 66884
rect 4876 66396 4940 66400
rect 4876 66340 4880 66396
rect 4880 66340 4936 66396
rect 4936 66340 4940 66396
rect 4876 66336 4940 66340
rect 4956 66396 5020 66400
rect 4956 66340 4960 66396
rect 4960 66340 5016 66396
rect 5016 66340 5020 66396
rect 4956 66336 5020 66340
rect 5036 66396 5100 66400
rect 5036 66340 5040 66396
rect 5040 66340 5096 66396
rect 5096 66340 5100 66396
rect 5036 66336 5100 66340
rect 5116 66396 5180 66400
rect 5116 66340 5120 66396
rect 5120 66340 5176 66396
rect 5176 66340 5180 66396
rect 5116 66336 5180 66340
rect 35596 66396 35660 66400
rect 35596 66340 35600 66396
rect 35600 66340 35656 66396
rect 35656 66340 35660 66396
rect 35596 66336 35660 66340
rect 35676 66396 35740 66400
rect 35676 66340 35680 66396
rect 35680 66340 35736 66396
rect 35736 66340 35740 66396
rect 35676 66336 35740 66340
rect 35756 66396 35820 66400
rect 35756 66340 35760 66396
rect 35760 66340 35816 66396
rect 35816 66340 35820 66396
rect 35756 66336 35820 66340
rect 35836 66396 35900 66400
rect 35836 66340 35840 66396
rect 35840 66340 35896 66396
rect 35896 66340 35900 66396
rect 35836 66336 35900 66340
rect 66316 66396 66380 66400
rect 66316 66340 66320 66396
rect 66320 66340 66376 66396
rect 66376 66340 66380 66396
rect 66316 66336 66380 66340
rect 66396 66396 66460 66400
rect 66396 66340 66400 66396
rect 66400 66340 66456 66396
rect 66456 66340 66460 66396
rect 66396 66336 66460 66340
rect 66476 66396 66540 66400
rect 66476 66340 66480 66396
rect 66480 66340 66536 66396
rect 66536 66340 66540 66396
rect 66476 66336 66540 66340
rect 66556 66396 66620 66400
rect 66556 66340 66560 66396
rect 66560 66340 66616 66396
rect 66616 66340 66620 66396
rect 66556 66336 66620 66340
rect 97036 66396 97100 66400
rect 97036 66340 97040 66396
rect 97040 66340 97096 66396
rect 97096 66340 97100 66396
rect 97036 66336 97100 66340
rect 97116 66396 97180 66400
rect 97116 66340 97120 66396
rect 97120 66340 97176 66396
rect 97176 66340 97180 66396
rect 97116 66336 97180 66340
rect 97196 66396 97260 66400
rect 97196 66340 97200 66396
rect 97200 66340 97256 66396
rect 97256 66340 97260 66396
rect 97196 66336 97260 66340
rect 97276 66396 97340 66400
rect 97276 66340 97280 66396
rect 97280 66340 97336 66396
rect 97336 66340 97340 66396
rect 97276 66336 97340 66340
rect 4216 65852 4280 65856
rect 4216 65796 4220 65852
rect 4220 65796 4276 65852
rect 4276 65796 4280 65852
rect 4216 65792 4280 65796
rect 4296 65852 4360 65856
rect 4296 65796 4300 65852
rect 4300 65796 4356 65852
rect 4356 65796 4360 65852
rect 4296 65792 4360 65796
rect 4376 65852 4440 65856
rect 4376 65796 4380 65852
rect 4380 65796 4436 65852
rect 4436 65796 4440 65852
rect 4376 65792 4440 65796
rect 4456 65852 4520 65856
rect 4456 65796 4460 65852
rect 4460 65796 4516 65852
rect 4516 65796 4520 65852
rect 4456 65792 4520 65796
rect 34936 65852 35000 65856
rect 34936 65796 34940 65852
rect 34940 65796 34996 65852
rect 34996 65796 35000 65852
rect 34936 65792 35000 65796
rect 35016 65852 35080 65856
rect 35016 65796 35020 65852
rect 35020 65796 35076 65852
rect 35076 65796 35080 65852
rect 35016 65792 35080 65796
rect 35096 65852 35160 65856
rect 35096 65796 35100 65852
rect 35100 65796 35156 65852
rect 35156 65796 35160 65852
rect 35096 65792 35160 65796
rect 35176 65852 35240 65856
rect 35176 65796 35180 65852
rect 35180 65796 35236 65852
rect 35236 65796 35240 65852
rect 35176 65792 35240 65796
rect 65656 65852 65720 65856
rect 65656 65796 65660 65852
rect 65660 65796 65716 65852
rect 65716 65796 65720 65852
rect 65656 65792 65720 65796
rect 65736 65852 65800 65856
rect 65736 65796 65740 65852
rect 65740 65796 65796 65852
rect 65796 65796 65800 65852
rect 65736 65792 65800 65796
rect 65816 65852 65880 65856
rect 65816 65796 65820 65852
rect 65820 65796 65876 65852
rect 65876 65796 65880 65852
rect 65816 65792 65880 65796
rect 65896 65852 65960 65856
rect 65896 65796 65900 65852
rect 65900 65796 65956 65852
rect 65956 65796 65960 65852
rect 65896 65792 65960 65796
rect 96376 65852 96440 65856
rect 96376 65796 96380 65852
rect 96380 65796 96436 65852
rect 96436 65796 96440 65852
rect 96376 65792 96440 65796
rect 96456 65852 96520 65856
rect 96456 65796 96460 65852
rect 96460 65796 96516 65852
rect 96516 65796 96520 65852
rect 96456 65792 96520 65796
rect 96536 65852 96600 65856
rect 96536 65796 96540 65852
rect 96540 65796 96596 65852
rect 96596 65796 96600 65852
rect 96536 65792 96600 65796
rect 96616 65852 96680 65856
rect 96616 65796 96620 65852
rect 96620 65796 96676 65852
rect 96676 65796 96680 65852
rect 96616 65792 96680 65796
rect 4876 65308 4940 65312
rect 4876 65252 4880 65308
rect 4880 65252 4936 65308
rect 4936 65252 4940 65308
rect 4876 65248 4940 65252
rect 4956 65308 5020 65312
rect 4956 65252 4960 65308
rect 4960 65252 5016 65308
rect 5016 65252 5020 65308
rect 4956 65248 5020 65252
rect 5036 65308 5100 65312
rect 5036 65252 5040 65308
rect 5040 65252 5096 65308
rect 5096 65252 5100 65308
rect 5036 65248 5100 65252
rect 5116 65308 5180 65312
rect 5116 65252 5120 65308
rect 5120 65252 5176 65308
rect 5176 65252 5180 65308
rect 5116 65248 5180 65252
rect 35596 65308 35660 65312
rect 35596 65252 35600 65308
rect 35600 65252 35656 65308
rect 35656 65252 35660 65308
rect 35596 65248 35660 65252
rect 35676 65308 35740 65312
rect 35676 65252 35680 65308
rect 35680 65252 35736 65308
rect 35736 65252 35740 65308
rect 35676 65248 35740 65252
rect 35756 65308 35820 65312
rect 35756 65252 35760 65308
rect 35760 65252 35816 65308
rect 35816 65252 35820 65308
rect 35756 65248 35820 65252
rect 35836 65308 35900 65312
rect 35836 65252 35840 65308
rect 35840 65252 35896 65308
rect 35896 65252 35900 65308
rect 35836 65248 35900 65252
rect 66316 65308 66380 65312
rect 66316 65252 66320 65308
rect 66320 65252 66376 65308
rect 66376 65252 66380 65308
rect 66316 65248 66380 65252
rect 66396 65308 66460 65312
rect 66396 65252 66400 65308
rect 66400 65252 66456 65308
rect 66456 65252 66460 65308
rect 66396 65248 66460 65252
rect 66476 65308 66540 65312
rect 66476 65252 66480 65308
rect 66480 65252 66536 65308
rect 66536 65252 66540 65308
rect 66476 65248 66540 65252
rect 66556 65308 66620 65312
rect 66556 65252 66560 65308
rect 66560 65252 66616 65308
rect 66616 65252 66620 65308
rect 66556 65248 66620 65252
rect 97036 65308 97100 65312
rect 97036 65252 97040 65308
rect 97040 65252 97096 65308
rect 97096 65252 97100 65308
rect 97036 65248 97100 65252
rect 97116 65308 97180 65312
rect 97116 65252 97120 65308
rect 97120 65252 97176 65308
rect 97176 65252 97180 65308
rect 97116 65248 97180 65252
rect 97196 65308 97260 65312
rect 97196 65252 97200 65308
rect 97200 65252 97256 65308
rect 97256 65252 97260 65308
rect 97196 65248 97260 65252
rect 97276 65308 97340 65312
rect 97276 65252 97280 65308
rect 97280 65252 97336 65308
rect 97336 65252 97340 65308
rect 97276 65248 97340 65252
rect 4216 64764 4280 64768
rect 4216 64708 4220 64764
rect 4220 64708 4276 64764
rect 4276 64708 4280 64764
rect 4216 64704 4280 64708
rect 4296 64764 4360 64768
rect 4296 64708 4300 64764
rect 4300 64708 4356 64764
rect 4356 64708 4360 64764
rect 4296 64704 4360 64708
rect 4376 64764 4440 64768
rect 4376 64708 4380 64764
rect 4380 64708 4436 64764
rect 4436 64708 4440 64764
rect 4376 64704 4440 64708
rect 4456 64764 4520 64768
rect 4456 64708 4460 64764
rect 4460 64708 4516 64764
rect 4516 64708 4520 64764
rect 4456 64704 4520 64708
rect 34936 64764 35000 64768
rect 34936 64708 34940 64764
rect 34940 64708 34996 64764
rect 34996 64708 35000 64764
rect 34936 64704 35000 64708
rect 35016 64764 35080 64768
rect 35016 64708 35020 64764
rect 35020 64708 35076 64764
rect 35076 64708 35080 64764
rect 35016 64704 35080 64708
rect 35096 64764 35160 64768
rect 35096 64708 35100 64764
rect 35100 64708 35156 64764
rect 35156 64708 35160 64764
rect 35096 64704 35160 64708
rect 35176 64764 35240 64768
rect 35176 64708 35180 64764
rect 35180 64708 35236 64764
rect 35236 64708 35240 64764
rect 35176 64704 35240 64708
rect 65656 64764 65720 64768
rect 65656 64708 65660 64764
rect 65660 64708 65716 64764
rect 65716 64708 65720 64764
rect 65656 64704 65720 64708
rect 65736 64764 65800 64768
rect 65736 64708 65740 64764
rect 65740 64708 65796 64764
rect 65796 64708 65800 64764
rect 65736 64704 65800 64708
rect 65816 64764 65880 64768
rect 65816 64708 65820 64764
rect 65820 64708 65876 64764
rect 65876 64708 65880 64764
rect 65816 64704 65880 64708
rect 65896 64764 65960 64768
rect 65896 64708 65900 64764
rect 65900 64708 65956 64764
rect 65956 64708 65960 64764
rect 65896 64704 65960 64708
rect 96376 64764 96440 64768
rect 96376 64708 96380 64764
rect 96380 64708 96436 64764
rect 96436 64708 96440 64764
rect 96376 64704 96440 64708
rect 96456 64764 96520 64768
rect 96456 64708 96460 64764
rect 96460 64708 96516 64764
rect 96516 64708 96520 64764
rect 96456 64704 96520 64708
rect 96536 64764 96600 64768
rect 96536 64708 96540 64764
rect 96540 64708 96596 64764
rect 96596 64708 96600 64764
rect 96536 64704 96600 64708
rect 96616 64764 96680 64768
rect 96616 64708 96620 64764
rect 96620 64708 96676 64764
rect 96676 64708 96680 64764
rect 96616 64704 96680 64708
rect 4876 64220 4940 64224
rect 4876 64164 4880 64220
rect 4880 64164 4936 64220
rect 4936 64164 4940 64220
rect 4876 64160 4940 64164
rect 4956 64220 5020 64224
rect 4956 64164 4960 64220
rect 4960 64164 5016 64220
rect 5016 64164 5020 64220
rect 4956 64160 5020 64164
rect 5036 64220 5100 64224
rect 5036 64164 5040 64220
rect 5040 64164 5096 64220
rect 5096 64164 5100 64220
rect 5036 64160 5100 64164
rect 5116 64220 5180 64224
rect 5116 64164 5120 64220
rect 5120 64164 5176 64220
rect 5176 64164 5180 64220
rect 5116 64160 5180 64164
rect 35596 64220 35660 64224
rect 35596 64164 35600 64220
rect 35600 64164 35656 64220
rect 35656 64164 35660 64220
rect 35596 64160 35660 64164
rect 35676 64220 35740 64224
rect 35676 64164 35680 64220
rect 35680 64164 35736 64220
rect 35736 64164 35740 64220
rect 35676 64160 35740 64164
rect 35756 64220 35820 64224
rect 35756 64164 35760 64220
rect 35760 64164 35816 64220
rect 35816 64164 35820 64220
rect 35756 64160 35820 64164
rect 35836 64220 35900 64224
rect 35836 64164 35840 64220
rect 35840 64164 35896 64220
rect 35896 64164 35900 64220
rect 35836 64160 35900 64164
rect 66316 64220 66380 64224
rect 66316 64164 66320 64220
rect 66320 64164 66376 64220
rect 66376 64164 66380 64220
rect 66316 64160 66380 64164
rect 66396 64220 66460 64224
rect 66396 64164 66400 64220
rect 66400 64164 66456 64220
rect 66456 64164 66460 64220
rect 66396 64160 66460 64164
rect 66476 64220 66540 64224
rect 66476 64164 66480 64220
rect 66480 64164 66536 64220
rect 66536 64164 66540 64220
rect 66476 64160 66540 64164
rect 66556 64220 66620 64224
rect 66556 64164 66560 64220
rect 66560 64164 66616 64220
rect 66616 64164 66620 64220
rect 66556 64160 66620 64164
rect 97036 64220 97100 64224
rect 97036 64164 97040 64220
rect 97040 64164 97096 64220
rect 97096 64164 97100 64220
rect 97036 64160 97100 64164
rect 97116 64220 97180 64224
rect 97116 64164 97120 64220
rect 97120 64164 97176 64220
rect 97176 64164 97180 64220
rect 97116 64160 97180 64164
rect 97196 64220 97260 64224
rect 97196 64164 97200 64220
rect 97200 64164 97256 64220
rect 97256 64164 97260 64220
rect 97196 64160 97260 64164
rect 97276 64220 97340 64224
rect 97276 64164 97280 64220
rect 97280 64164 97336 64220
rect 97336 64164 97340 64220
rect 97276 64160 97340 64164
rect 4216 63676 4280 63680
rect 4216 63620 4220 63676
rect 4220 63620 4276 63676
rect 4276 63620 4280 63676
rect 4216 63616 4280 63620
rect 4296 63676 4360 63680
rect 4296 63620 4300 63676
rect 4300 63620 4356 63676
rect 4356 63620 4360 63676
rect 4296 63616 4360 63620
rect 4376 63676 4440 63680
rect 4376 63620 4380 63676
rect 4380 63620 4436 63676
rect 4436 63620 4440 63676
rect 4376 63616 4440 63620
rect 4456 63676 4520 63680
rect 4456 63620 4460 63676
rect 4460 63620 4516 63676
rect 4516 63620 4520 63676
rect 4456 63616 4520 63620
rect 34936 63676 35000 63680
rect 34936 63620 34940 63676
rect 34940 63620 34996 63676
rect 34996 63620 35000 63676
rect 34936 63616 35000 63620
rect 35016 63676 35080 63680
rect 35016 63620 35020 63676
rect 35020 63620 35076 63676
rect 35076 63620 35080 63676
rect 35016 63616 35080 63620
rect 35096 63676 35160 63680
rect 35096 63620 35100 63676
rect 35100 63620 35156 63676
rect 35156 63620 35160 63676
rect 35096 63616 35160 63620
rect 35176 63676 35240 63680
rect 35176 63620 35180 63676
rect 35180 63620 35236 63676
rect 35236 63620 35240 63676
rect 35176 63616 35240 63620
rect 65656 63676 65720 63680
rect 65656 63620 65660 63676
rect 65660 63620 65716 63676
rect 65716 63620 65720 63676
rect 65656 63616 65720 63620
rect 65736 63676 65800 63680
rect 65736 63620 65740 63676
rect 65740 63620 65796 63676
rect 65796 63620 65800 63676
rect 65736 63616 65800 63620
rect 65816 63676 65880 63680
rect 65816 63620 65820 63676
rect 65820 63620 65876 63676
rect 65876 63620 65880 63676
rect 65816 63616 65880 63620
rect 65896 63676 65960 63680
rect 65896 63620 65900 63676
rect 65900 63620 65956 63676
rect 65956 63620 65960 63676
rect 65896 63616 65960 63620
rect 96376 63676 96440 63680
rect 96376 63620 96380 63676
rect 96380 63620 96436 63676
rect 96436 63620 96440 63676
rect 96376 63616 96440 63620
rect 96456 63676 96520 63680
rect 96456 63620 96460 63676
rect 96460 63620 96516 63676
rect 96516 63620 96520 63676
rect 96456 63616 96520 63620
rect 96536 63676 96600 63680
rect 96536 63620 96540 63676
rect 96540 63620 96596 63676
rect 96596 63620 96600 63676
rect 96536 63616 96600 63620
rect 96616 63676 96680 63680
rect 96616 63620 96620 63676
rect 96620 63620 96676 63676
rect 96676 63620 96680 63676
rect 96616 63616 96680 63620
rect 4876 63132 4940 63136
rect 4876 63076 4880 63132
rect 4880 63076 4936 63132
rect 4936 63076 4940 63132
rect 4876 63072 4940 63076
rect 4956 63132 5020 63136
rect 4956 63076 4960 63132
rect 4960 63076 5016 63132
rect 5016 63076 5020 63132
rect 4956 63072 5020 63076
rect 5036 63132 5100 63136
rect 5036 63076 5040 63132
rect 5040 63076 5096 63132
rect 5096 63076 5100 63132
rect 5036 63072 5100 63076
rect 5116 63132 5180 63136
rect 5116 63076 5120 63132
rect 5120 63076 5176 63132
rect 5176 63076 5180 63132
rect 5116 63072 5180 63076
rect 35596 63132 35660 63136
rect 35596 63076 35600 63132
rect 35600 63076 35656 63132
rect 35656 63076 35660 63132
rect 35596 63072 35660 63076
rect 35676 63132 35740 63136
rect 35676 63076 35680 63132
rect 35680 63076 35736 63132
rect 35736 63076 35740 63132
rect 35676 63072 35740 63076
rect 35756 63132 35820 63136
rect 35756 63076 35760 63132
rect 35760 63076 35816 63132
rect 35816 63076 35820 63132
rect 35756 63072 35820 63076
rect 35836 63132 35900 63136
rect 35836 63076 35840 63132
rect 35840 63076 35896 63132
rect 35896 63076 35900 63132
rect 35836 63072 35900 63076
rect 66316 63132 66380 63136
rect 66316 63076 66320 63132
rect 66320 63076 66376 63132
rect 66376 63076 66380 63132
rect 66316 63072 66380 63076
rect 66396 63132 66460 63136
rect 66396 63076 66400 63132
rect 66400 63076 66456 63132
rect 66456 63076 66460 63132
rect 66396 63072 66460 63076
rect 66476 63132 66540 63136
rect 66476 63076 66480 63132
rect 66480 63076 66536 63132
rect 66536 63076 66540 63132
rect 66476 63072 66540 63076
rect 66556 63132 66620 63136
rect 66556 63076 66560 63132
rect 66560 63076 66616 63132
rect 66616 63076 66620 63132
rect 66556 63072 66620 63076
rect 97036 63132 97100 63136
rect 97036 63076 97040 63132
rect 97040 63076 97096 63132
rect 97096 63076 97100 63132
rect 97036 63072 97100 63076
rect 97116 63132 97180 63136
rect 97116 63076 97120 63132
rect 97120 63076 97176 63132
rect 97176 63076 97180 63132
rect 97116 63072 97180 63076
rect 97196 63132 97260 63136
rect 97196 63076 97200 63132
rect 97200 63076 97256 63132
rect 97256 63076 97260 63132
rect 97196 63072 97260 63076
rect 97276 63132 97340 63136
rect 97276 63076 97280 63132
rect 97280 63076 97336 63132
rect 97336 63076 97340 63132
rect 97276 63072 97340 63076
rect 35388 62732 35452 62796
rect 4216 62588 4280 62592
rect 4216 62532 4220 62588
rect 4220 62532 4276 62588
rect 4276 62532 4280 62588
rect 4216 62528 4280 62532
rect 4296 62588 4360 62592
rect 4296 62532 4300 62588
rect 4300 62532 4356 62588
rect 4356 62532 4360 62588
rect 4296 62528 4360 62532
rect 4376 62588 4440 62592
rect 4376 62532 4380 62588
rect 4380 62532 4436 62588
rect 4436 62532 4440 62588
rect 4376 62528 4440 62532
rect 4456 62588 4520 62592
rect 4456 62532 4460 62588
rect 4460 62532 4516 62588
rect 4516 62532 4520 62588
rect 4456 62528 4520 62532
rect 34936 62588 35000 62592
rect 34936 62532 34940 62588
rect 34940 62532 34996 62588
rect 34996 62532 35000 62588
rect 34936 62528 35000 62532
rect 35016 62588 35080 62592
rect 35016 62532 35020 62588
rect 35020 62532 35076 62588
rect 35076 62532 35080 62588
rect 35016 62528 35080 62532
rect 35096 62588 35160 62592
rect 35096 62532 35100 62588
rect 35100 62532 35156 62588
rect 35156 62532 35160 62588
rect 35096 62528 35160 62532
rect 35176 62588 35240 62592
rect 35176 62532 35180 62588
rect 35180 62532 35236 62588
rect 35236 62532 35240 62588
rect 35176 62528 35240 62532
rect 65656 62588 65720 62592
rect 65656 62532 65660 62588
rect 65660 62532 65716 62588
rect 65716 62532 65720 62588
rect 65656 62528 65720 62532
rect 65736 62588 65800 62592
rect 65736 62532 65740 62588
rect 65740 62532 65796 62588
rect 65796 62532 65800 62588
rect 65736 62528 65800 62532
rect 65816 62588 65880 62592
rect 65816 62532 65820 62588
rect 65820 62532 65876 62588
rect 65876 62532 65880 62588
rect 65816 62528 65880 62532
rect 65896 62588 65960 62592
rect 65896 62532 65900 62588
rect 65900 62532 65956 62588
rect 65956 62532 65960 62588
rect 65896 62528 65960 62532
rect 96376 62588 96440 62592
rect 96376 62532 96380 62588
rect 96380 62532 96436 62588
rect 96436 62532 96440 62588
rect 96376 62528 96440 62532
rect 96456 62588 96520 62592
rect 96456 62532 96460 62588
rect 96460 62532 96516 62588
rect 96516 62532 96520 62588
rect 96456 62528 96520 62532
rect 96536 62588 96600 62592
rect 96536 62532 96540 62588
rect 96540 62532 96596 62588
rect 96596 62532 96600 62588
rect 96536 62528 96600 62532
rect 96616 62588 96680 62592
rect 96616 62532 96620 62588
rect 96620 62532 96676 62588
rect 96676 62532 96680 62588
rect 96616 62528 96680 62532
rect 4876 62044 4940 62048
rect 4876 61988 4880 62044
rect 4880 61988 4936 62044
rect 4936 61988 4940 62044
rect 4876 61984 4940 61988
rect 4956 62044 5020 62048
rect 4956 61988 4960 62044
rect 4960 61988 5016 62044
rect 5016 61988 5020 62044
rect 4956 61984 5020 61988
rect 5036 62044 5100 62048
rect 5036 61988 5040 62044
rect 5040 61988 5096 62044
rect 5096 61988 5100 62044
rect 5036 61984 5100 61988
rect 5116 62044 5180 62048
rect 5116 61988 5120 62044
rect 5120 61988 5176 62044
rect 5176 61988 5180 62044
rect 5116 61984 5180 61988
rect 35596 62044 35660 62048
rect 35596 61988 35600 62044
rect 35600 61988 35656 62044
rect 35656 61988 35660 62044
rect 35596 61984 35660 61988
rect 35676 62044 35740 62048
rect 35676 61988 35680 62044
rect 35680 61988 35736 62044
rect 35736 61988 35740 62044
rect 35676 61984 35740 61988
rect 35756 62044 35820 62048
rect 35756 61988 35760 62044
rect 35760 61988 35816 62044
rect 35816 61988 35820 62044
rect 35756 61984 35820 61988
rect 35836 62044 35900 62048
rect 35836 61988 35840 62044
rect 35840 61988 35896 62044
rect 35896 61988 35900 62044
rect 35836 61984 35900 61988
rect 66316 62044 66380 62048
rect 66316 61988 66320 62044
rect 66320 61988 66376 62044
rect 66376 61988 66380 62044
rect 66316 61984 66380 61988
rect 66396 62044 66460 62048
rect 66396 61988 66400 62044
rect 66400 61988 66456 62044
rect 66456 61988 66460 62044
rect 66396 61984 66460 61988
rect 66476 62044 66540 62048
rect 66476 61988 66480 62044
rect 66480 61988 66536 62044
rect 66536 61988 66540 62044
rect 66476 61984 66540 61988
rect 66556 62044 66620 62048
rect 66556 61988 66560 62044
rect 66560 61988 66616 62044
rect 66616 61988 66620 62044
rect 66556 61984 66620 61988
rect 97036 62044 97100 62048
rect 97036 61988 97040 62044
rect 97040 61988 97096 62044
rect 97096 61988 97100 62044
rect 97036 61984 97100 61988
rect 97116 62044 97180 62048
rect 97116 61988 97120 62044
rect 97120 61988 97176 62044
rect 97176 61988 97180 62044
rect 97116 61984 97180 61988
rect 97196 62044 97260 62048
rect 97196 61988 97200 62044
rect 97200 61988 97256 62044
rect 97256 61988 97260 62044
rect 97196 61984 97260 61988
rect 97276 62044 97340 62048
rect 97276 61988 97280 62044
rect 97280 61988 97336 62044
rect 97336 61988 97340 62044
rect 97276 61984 97340 61988
rect 4216 61500 4280 61504
rect 4216 61444 4220 61500
rect 4220 61444 4276 61500
rect 4276 61444 4280 61500
rect 4216 61440 4280 61444
rect 4296 61500 4360 61504
rect 4296 61444 4300 61500
rect 4300 61444 4356 61500
rect 4356 61444 4360 61500
rect 4296 61440 4360 61444
rect 4376 61500 4440 61504
rect 4376 61444 4380 61500
rect 4380 61444 4436 61500
rect 4436 61444 4440 61500
rect 4376 61440 4440 61444
rect 4456 61500 4520 61504
rect 4456 61444 4460 61500
rect 4460 61444 4516 61500
rect 4516 61444 4520 61500
rect 4456 61440 4520 61444
rect 34936 61500 35000 61504
rect 34936 61444 34940 61500
rect 34940 61444 34996 61500
rect 34996 61444 35000 61500
rect 34936 61440 35000 61444
rect 35016 61500 35080 61504
rect 35016 61444 35020 61500
rect 35020 61444 35076 61500
rect 35076 61444 35080 61500
rect 35016 61440 35080 61444
rect 35096 61500 35160 61504
rect 35096 61444 35100 61500
rect 35100 61444 35156 61500
rect 35156 61444 35160 61500
rect 35096 61440 35160 61444
rect 35176 61500 35240 61504
rect 35176 61444 35180 61500
rect 35180 61444 35236 61500
rect 35236 61444 35240 61500
rect 35176 61440 35240 61444
rect 65656 61500 65720 61504
rect 65656 61444 65660 61500
rect 65660 61444 65716 61500
rect 65716 61444 65720 61500
rect 65656 61440 65720 61444
rect 65736 61500 65800 61504
rect 65736 61444 65740 61500
rect 65740 61444 65796 61500
rect 65796 61444 65800 61500
rect 65736 61440 65800 61444
rect 65816 61500 65880 61504
rect 65816 61444 65820 61500
rect 65820 61444 65876 61500
rect 65876 61444 65880 61500
rect 65816 61440 65880 61444
rect 65896 61500 65960 61504
rect 65896 61444 65900 61500
rect 65900 61444 65956 61500
rect 65956 61444 65960 61500
rect 65896 61440 65960 61444
rect 96376 61500 96440 61504
rect 96376 61444 96380 61500
rect 96380 61444 96436 61500
rect 96436 61444 96440 61500
rect 96376 61440 96440 61444
rect 96456 61500 96520 61504
rect 96456 61444 96460 61500
rect 96460 61444 96516 61500
rect 96516 61444 96520 61500
rect 96456 61440 96520 61444
rect 96536 61500 96600 61504
rect 96536 61444 96540 61500
rect 96540 61444 96596 61500
rect 96596 61444 96600 61500
rect 96536 61440 96600 61444
rect 96616 61500 96680 61504
rect 96616 61444 96620 61500
rect 96620 61444 96676 61500
rect 96676 61444 96680 61500
rect 96616 61440 96680 61444
rect 4876 60956 4940 60960
rect 4876 60900 4880 60956
rect 4880 60900 4936 60956
rect 4936 60900 4940 60956
rect 4876 60896 4940 60900
rect 4956 60956 5020 60960
rect 4956 60900 4960 60956
rect 4960 60900 5016 60956
rect 5016 60900 5020 60956
rect 4956 60896 5020 60900
rect 5036 60956 5100 60960
rect 5036 60900 5040 60956
rect 5040 60900 5096 60956
rect 5096 60900 5100 60956
rect 5036 60896 5100 60900
rect 5116 60956 5180 60960
rect 5116 60900 5120 60956
rect 5120 60900 5176 60956
rect 5176 60900 5180 60956
rect 5116 60896 5180 60900
rect 35596 60956 35660 60960
rect 35596 60900 35600 60956
rect 35600 60900 35656 60956
rect 35656 60900 35660 60956
rect 35596 60896 35660 60900
rect 35676 60956 35740 60960
rect 35676 60900 35680 60956
rect 35680 60900 35736 60956
rect 35736 60900 35740 60956
rect 35676 60896 35740 60900
rect 35756 60956 35820 60960
rect 35756 60900 35760 60956
rect 35760 60900 35816 60956
rect 35816 60900 35820 60956
rect 35756 60896 35820 60900
rect 35836 60956 35900 60960
rect 35836 60900 35840 60956
rect 35840 60900 35896 60956
rect 35896 60900 35900 60956
rect 35836 60896 35900 60900
rect 66316 60956 66380 60960
rect 66316 60900 66320 60956
rect 66320 60900 66376 60956
rect 66376 60900 66380 60956
rect 66316 60896 66380 60900
rect 66396 60956 66460 60960
rect 66396 60900 66400 60956
rect 66400 60900 66456 60956
rect 66456 60900 66460 60956
rect 66396 60896 66460 60900
rect 66476 60956 66540 60960
rect 66476 60900 66480 60956
rect 66480 60900 66536 60956
rect 66536 60900 66540 60956
rect 66476 60896 66540 60900
rect 66556 60956 66620 60960
rect 66556 60900 66560 60956
rect 66560 60900 66616 60956
rect 66616 60900 66620 60956
rect 66556 60896 66620 60900
rect 97036 60956 97100 60960
rect 97036 60900 97040 60956
rect 97040 60900 97096 60956
rect 97096 60900 97100 60956
rect 97036 60896 97100 60900
rect 97116 60956 97180 60960
rect 97116 60900 97120 60956
rect 97120 60900 97176 60956
rect 97176 60900 97180 60956
rect 97116 60896 97180 60900
rect 97196 60956 97260 60960
rect 97196 60900 97200 60956
rect 97200 60900 97256 60956
rect 97256 60900 97260 60956
rect 97196 60896 97260 60900
rect 97276 60956 97340 60960
rect 97276 60900 97280 60956
rect 97280 60900 97336 60956
rect 97336 60900 97340 60956
rect 97276 60896 97340 60900
rect 67588 60692 67652 60756
rect 1308 60412 1372 60416
rect 1308 60356 1312 60412
rect 1312 60356 1368 60412
rect 1368 60356 1372 60412
rect 1308 60352 1372 60356
rect 1388 60412 1452 60416
rect 1388 60356 1392 60412
rect 1392 60356 1448 60412
rect 1448 60356 1452 60412
rect 1388 60352 1452 60356
rect 4216 60412 4280 60416
rect 4216 60356 4220 60412
rect 4220 60356 4276 60412
rect 4276 60356 4280 60412
rect 4216 60352 4280 60356
rect 4296 60412 4360 60416
rect 4296 60356 4300 60412
rect 4300 60356 4356 60412
rect 4356 60356 4360 60412
rect 4296 60352 4360 60356
rect 4376 60412 4440 60416
rect 4376 60356 4380 60412
rect 4380 60356 4436 60412
rect 4436 60356 4440 60412
rect 4376 60352 4440 60356
rect 4456 60412 4520 60416
rect 4456 60356 4460 60412
rect 4460 60356 4516 60412
rect 4516 60356 4520 60412
rect 4456 60352 4520 60356
rect 34936 60412 35000 60416
rect 34936 60356 34940 60412
rect 34940 60356 34996 60412
rect 34996 60356 35000 60412
rect 34936 60352 35000 60356
rect 35016 60412 35080 60416
rect 35016 60356 35020 60412
rect 35020 60356 35076 60412
rect 35076 60356 35080 60412
rect 35016 60352 35080 60356
rect 35096 60412 35160 60416
rect 35096 60356 35100 60412
rect 35100 60356 35156 60412
rect 35156 60356 35160 60412
rect 35096 60352 35160 60356
rect 35176 60412 35240 60416
rect 35176 60356 35180 60412
rect 35180 60356 35236 60412
rect 35236 60356 35240 60412
rect 35176 60352 35240 60356
rect 65656 60412 65720 60416
rect 65656 60356 65660 60412
rect 65660 60356 65716 60412
rect 65716 60356 65720 60412
rect 65656 60352 65720 60356
rect 65736 60412 65800 60416
rect 65736 60356 65740 60412
rect 65740 60356 65796 60412
rect 65796 60356 65800 60412
rect 65736 60352 65800 60356
rect 65816 60412 65880 60416
rect 65816 60356 65820 60412
rect 65820 60356 65876 60412
rect 65876 60356 65880 60412
rect 65816 60352 65880 60356
rect 65896 60412 65960 60416
rect 65896 60356 65900 60412
rect 65900 60356 65956 60412
rect 65956 60356 65960 60412
rect 65896 60352 65960 60356
rect 96376 60412 96440 60416
rect 96376 60356 96380 60412
rect 96380 60356 96436 60412
rect 96436 60356 96440 60412
rect 96376 60352 96440 60356
rect 96456 60412 96520 60416
rect 96456 60356 96460 60412
rect 96460 60356 96516 60412
rect 96516 60356 96520 60412
rect 96456 60352 96520 60356
rect 96536 60412 96600 60416
rect 96536 60356 96540 60412
rect 96540 60356 96596 60412
rect 96596 60356 96600 60412
rect 96536 60352 96600 60356
rect 96616 60412 96680 60416
rect 96616 60356 96620 60412
rect 96620 60356 96676 60412
rect 96676 60356 96680 60412
rect 96616 60352 96680 60356
rect 98932 60412 98996 60416
rect 98932 60356 98936 60412
rect 98936 60356 98992 60412
rect 98992 60356 98996 60412
rect 98932 60352 98996 60356
rect 99012 60412 99076 60416
rect 99012 60356 99016 60412
rect 99016 60356 99072 60412
rect 99072 60356 99076 60412
rect 99012 60352 99076 60356
rect 99092 60412 99156 60416
rect 99092 60356 99096 60412
rect 99096 60356 99152 60412
rect 99152 60356 99156 60412
rect 99092 60352 99156 60356
rect 99172 60412 99236 60416
rect 99172 60356 99176 60412
rect 99176 60356 99232 60412
rect 99232 60356 99236 60412
rect 99172 60352 99236 60356
rect 1676 59868 1740 59872
rect 1676 59812 1680 59868
rect 1680 59812 1736 59868
rect 1736 59812 1740 59868
rect 1676 59808 1740 59812
rect 1756 59868 1820 59872
rect 1756 59812 1760 59868
rect 1760 59812 1816 59868
rect 1816 59812 1820 59868
rect 1756 59808 1820 59812
rect 4876 59868 4940 59872
rect 4876 59812 4880 59868
rect 4880 59812 4936 59868
rect 4936 59812 4940 59868
rect 4876 59808 4940 59812
rect 4956 59868 5020 59872
rect 4956 59812 4960 59868
rect 4960 59812 5016 59868
rect 5016 59812 5020 59868
rect 4956 59808 5020 59812
rect 5036 59868 5100 59872
rect 5036 59812 5040 59868
rect 5040 59812 5096 59868
rect 5096 59812 5100 59868
rect 5036 59808 5100 59812
rect 5116 59868 5180 59872
rect 5116 59812 5120 59868
rect 5120 59812 5176 59868
rect 5176 59812 5180 59868
rect 5116 59808 5180 59812
rect 35596 59868 35660 59872
rect 35596 59812 35600 59868
rect 35600 59812 35656 59868
rect 35656 59812 35660 59868
rect 35596 59808 35660 59812
rect 35676 59868 35740 59872
rect 35676 59812 35680 59868
rect 35680 59812 35736 59868
rect 35736 59812 35740 59868
rect 35676 59808 35740 59812
rect 35756 59868 35820 59872
rect 35756 59812 35760 59868
rect 35760 59812 35816 59868
rect 35816 59812 35820 59868
rect 35756 59808 35820 59812
rect 35836 59868 35900 59872
rect 35836 59812 35840 59868
rect 35840 59812 35896 59868
rect 35896 59812 35900 59868
rect 35836 59808 35900 59812
rect 66316 59868 66380 59872
rect 66316 59812 66320 59868
rect 66320 59812 66376 59868
rect 66376 59812 66380 59868
rect 66316 59808 66380 59812
rect 66396 59868 66460 59872
rect 66396 59812 66400 59868
rect 66400 59812 66456 59868
rect 66456 59812 66460 59868
rect 66396 59808 66460 59812
rect 66476 59868 66540 59872
rect 66476 59812 66480 59868
rect 66480 59812 66536 59868
rect 66536 59812 66540 59868
rect 66476 59808 66540 59812
rect 66556 59868 66620 59872
rect 66556 59812 66560 59868
rect 66560 59812 66616 59868
rect 66616 59812 66620 59868
rect 66556 59808 66620 59812
rect 97036 59868 97100 59872
rect 97036 59812 97040 59868
rect 97040 59812 97096 59868
rect 97096 59812 97100 59868
rect 97036 59808 97100 59812
rect 97116 59868 97180 59872
rect 97116 59812 97120 59868
rect 97120 59812 97176 59868
rect 97176 59812 97180 59868
rect 97116 59808 97180 59812
rect 97196 59868 97260 59872
rect 97196 59812 97200 59868
rect 97200 59812 97256 59868
rect 97256 59812 97260 59868
rect 97196 59808 97260 59812
rect 97276 59868 97340 59872
rect 97276 59812 97280 59868
rect 97280 59812 97336 59868
rect 97336 59812 97340 59868
rect 97276 59808 97340 59812
rect 99668 59868 99732 59872
rect 99668 59812 99672 59868
rect 99672 59812 99728 59868
rect 99728 59812 99732 59868
rect 99668 59808 99732 59812
rect 99748 59868 99812 59872
rect 99748 59812 99752 59868
rect 99752 59812 99808 59868
rect 99808 59812 99812 59868
rect 99748 59808 99812 59812
rect 99828 59868 99892 59872
rect 99828 59812 99832 59868
rect 99832 59812 99888 59868
rect 99888 59812 99892 59868
rect 99828 59808 99892 59812
rect 99908 59868 99972 59872
rect 99908 59812 99912 59868
rect 99912 59812 99968 59868
rect 99968 59812 99972 59868
rect 99908 59808 99972 59812
rect 1308 59324 1372 59328
rect 1308 59268 1312 59324
rect 1312 59268 1368 59324
rect 1368 59268 1372 59324
rect 1308 59264 1372 59268
rect 1388 59324 1452 59328
rect 1388 59268 1392 59324
rect 1392 59268 1448 59324
rect 1448 59268 1452 59324
rect 1388 59264 1452 59268
rect 98932 59324 98996 59328
rect 98932 59268 98936 59324
rect 98936 59268 98992 59324
rect 98992 59268 98996 59324
rect 98932 59264 98996 59268
rect 99012 59324 99076 59328
rect 99012 59268 99016 59324
rect 99016 59268 99072 59324
rect 99072 59268 99076 59324
rect 99012 59264 99076 59268
rect 99092 59324 99156 59328
rect 99092 59268 99096 59324
rect 99096 59268 99152 59324
rect 99152 59268 99156 59324
rect 99092 59264 99156 59268
rect 99172 59324 99236 59328
rect 99172 59268 99176 59324
rect 99176 59268 99232 59324
rect 99232 59268 99236 59324
rect 99172 59264 99236 59268
rect 57468 58788 57532 58852
rect 1676 58780 1740 58784
rect 1676 58724 1680 58780
rect 1680 58724 1736 58780
rect 1736 58724 1740 58780
rect 1676 58720 1740 58724
rect 1756 58780 1820 58784
rect 1756 58724 1760 58780
rect 1760 58724 1816 58780
rect 1816 58724 1820 58780
rect 1756 58720 1820 58724
rect 99668 58780 99732 58784
rect 99668 58724 99672 58780
rect 99672 58724 99728 58780
rect 99728 58724 99732 58780
rect 99668 58720 99732 58724
rect 99748 58780 99812 58784
rect 99748 58724 99752 58780
rect 99752 58724 99808 58780
rect 99808 58724 99812 58780
rect 99748 58720 99812 58724
rect 99828 58780 99892 58784
rect 99828 58724 99832 58780
rect 99832 58724 99888 58780
rect 99888 58724 99892 58780
rect 99828 58720 99892 58724
rect 99908 58780 99972 58784
rect 99908 58724 99912 58780
rect 99912 58724 99968 58780
rect 99968 58724 99972 58780
rect 99908 58720 99972 58724
rect 62620 58652 62684 58716
rect 60044 58516 60108 58580
rect 1308 58236 1372 58240
rect 1308 58180 1312 58236
rect 1312 58180 1368 58236
rect 1368 58180 1372 58236
rect 1308 58176 1372 58180
rect 1388 58236 1452 58240
rect 1388 58180 1392 58236
rect 1392 58180 1448 58236
rect 1448 58180 1452 58236
rect 1388 58176 1452 58180
rect 98932 58236 98996 58240
rect 98932 58180 98936 58236
rect 98936 58180 98992 58236
rect 98992 58180 98996 58236
rect 98932 58176 98996 58180
rect 99012 58236 99076 58240
rect 99012 58180 99016 58236
rect 99016 58180 99072 58236
rect 99072 58180 99076 58236
rect 99012 58176 99076 58180
rect 99092 58236 99156 58240
rect 99092 58180 99096 58236
rect 99096 58180 99152 58236
rect 99152 58180 99156 58236
rect 99092 58176 99156 58180
rect 99172 58236 99236 58240
rect 99172 58180 99176 58236
rect 99176 58180 99232 58236
rect 99232 58180 99236 58236
rect 99172 58176 99236 58180
rect 32571 58108 32635 58172
rect 80142 58108 80206 58172
rect 81310 57972 81374 58036
rect 30075 57836 30139 57900
rect 65019 57836 65083 57900
rect 89858 57836 89922 57900
rect 1676 57692 1740 57696
rect 1676 57636 1680 57692
rect 1680 57636 1736 57692
rect 1736 57636 1740 57692
rect 1676 57632 1740 57636
rect 1756 57692 1820 57696
rect 1756 57636 1760 57692
rect 1760 57636 1816 57692
rect 1816 57636 1820 57692
rect 1756 57632 1820 57636
rect 99668 57692 99732 57696
rect 99668 57636 99672 57692
rect 99672 57636 99728 57692
rect 99728 57636 99732 57692
rect 99668 57632 99732 57636
rect 99748 57692 99812 57696
rect 99748 57636 99752 57692
rect 99752 57636 99808 57692
rect 99808 57636 99812 57692
rect 99748 57632 99812 57636
rect 99828 57692 99892 57696
rect 99828 57636 99832 57692
rect 99832 57636 99888 57692
rect 99888 57636 99892 57692
rect 99828 57632 99892 57636
rect 99908 57692 99972 57696
rect 99908 57636 99912 57692
rect 99912 57636 99968 57692
rect 99968 57636 99972 57692
rect 99908 57632 99972 57636
rect 1308 57148 1372 57152
rect 1308 57092 1312 57148
rect 1312 57092 1368 57148
rect 1368 57092 1372 57148
rect 1308 57088 1372 57092
rect 1388 57148 1452 57152
rect 1388 57092 1392 57148
rect 1392 57092 1448 57148
rect 1448 57092 1452 57148
rect 1388 57088 1452 57092
rect 98932 57148 98996 57152
rect 98932 57092 98936 57148
rect 98936 57092 98992 57148
rect 98992 57092 98996 57148
rect 98932 57088 98996 57092
rect 99012 57148 99076 57152
rect 99012 57092 99016 57148
rect 99016 57092 99072 57148
rect 99072 57092 99076 57148
rect 99012 57088 99076 57092
rect 99092 57148 99156 57152
rect 99092 57092 99096 57148
rect 99096 57092 99152 57148
rect 99152 57092 99156 57148
rect 99092 57088 99156 57092
rect 99172 57148 99236 57152
rect 99172 57092 99176 57148
rect 99176 57092 99232 57148
rect 99232 57092 99236 57148
rect 99172 57088 99236 57092
rect 1676 56604 1740 56608
rect 1676 56548 1680 56604
rect 1680 56548 1736 56604
rect 1736 56548 1740 56604
rect 1676 56544 1740 56548
rect 1756 56604 1820 56608
rect 1756 56548 1760 56604
rect 1760 56548 1816 56604
rect 1816 56548 1820 56604
rect 1756 56544 1820 56548
rect 99668 56604 99732 56608
rect 99668 56548 99672 56604
rect 99672 56548 99728 56604
rect 99728 56548 99732 56604
rect 99668 56544 99732 56548
rect 99748 56604 99812 56608
rect 99748 56548 99752 56604
rect 99752 56548 99808 56604
rect 99808 56548 99812 56604
rect 99748 56544 99812 56548
rect 99828 56604 99892 56608
rect 99828 56548 99832 56604
rect 99832 56548 99888 56604
rect 99888 56548 99892 56604
rect 99828 56544 99892 56548
rect 99908 56604 99972 56608
rect 99908 56548 99912 56604
rect 99912 56548 99968 56604
rect 99968 56548 99972 56604
rect 99908 56544 99972 56548
rect 1308 56060 1372 56064
rect 1308 56004 1312 56060
rect 1312 56004 1368 56060
rect 1368 56004 1372 56060
rect 1308 56000 1372 56004
rect 1388 56060 1452 56064
rect 1388 56004 1392 56060
rect 1392 56004 1448 56060
rect 1448 56004 1452 56060
rect 1388 56000 1452 56004
rect 98932 56060 98996 56064
rect 98932 56004 98936 56060
rect 98936 56004 98992 56060
rect 98992 56004 98996 56060
rect 98932 56000 98996 56004
rect 99012 56060 99076 56064
rect 99012 56004 99016 56060
rect 99016 56004 99072 56060
rect 99072 56004 99076 56060
rect 99012 56000 99076 56004
rect 99092 56060 99156 56064
rect 99092 56004 99096 56060
rect 99096 56004 99152 56060
rect 99152 56004 99156 56060
rect 99092 56000 99156 56004
rect 99172 56060 99236 56064
rect 99172 56004 99176 56060
rect 99176 56004 99232 56060
rect 99232 56004 99236 56060
rect 99172 56000 99236 56004
rect 1676 55516 1740 55520
rect 1676 55460 1680 55516
rect 1680 55460 1736 55516
rect 1736 55460 1740 55516
rect 1676 55456 1740 55460
rect 1756 55516 1820 55520
rect 1756 55460 1760 55516
rect 1760 55460 1816 55516
rect 1816 55460 1820 55516
rect 1756 55456 1820 55460
rect 99668 55516 99732 55520
rect 99668 55460 99672 55516
rect 99672 55460 99728 55516
rect 99728 55460 99732 55516
rect 99668 55456 99732 55460
rect 99748 55516 99812 55520
rect 99748 55460 99752 55516
rect 99752 55460 99808 55516
rect 99808 55460 99812 55516
rect 99748 55456 99812 55460
rect 99828 55516 99892 55520
rect 99828 55460 99832 55516
rect 99832 55460 99888 55516
rect 99888 55460 99892 55516
rect 99828 55456 99892 55460
rect 99908 55516 99972 55520
rect 99908 55460 99912 55516
rect 99912 55460 99968 55516
rect 99968 55460 99972 55516
rect 99908 55456 99972 55460
rect 1308 54972 1372 54976
rect 1308 54916 1312 54972
rect 1312 54916 1368 54972
rect 1368 54916 1372 54972
rect 1308 54912 1372 54916
rect 1388 54972 1452 54976
rect 1388 54916 1392 54972
rect 1392 54916 1448 54972
rect 1448 54916 1452 54972
rect 1388 54912 1452 54916
rect 98932 54972 98996 54976
rect 98932 54916 98936 54972
rect 98936 54916 98992 54972
rect 98992 54916 98996 54972
rect 98932 54912 98996 54916
rect 99012 54972 99076 54976
rect 99012 54916 99016 54972
rect 99016 54916 99072 54972
rect 99072 54916 99076 54972
rect 99012 54912 99076 54916
rect 99092 54972 99156 54976
rect 99092 54916 99096 54972
rect 99096 54916 99152 54972
rect 99152 54916 99156 54972
rect 99092 54912 99156 54916
rect 99172 54972 99236 54976
rect 99172 54916 99176 54972
rect 99176 54916 99232 54972
rect 99232 54916 99236 54972
rect 99172 54912 99236 54916
rect 1676 54428 1740 54432
rect 1676 54372 1680 54428
rect 1680 54372 1736 54428
rect 1736 54372 1740 54428
rect 1676 54368 1740 54372
rect 1756 54428 1820 54432
rect 1756 54372 1760 54428
rect 1760 54372 1816 54428
rect 1816 54372 1820 54428
rect 1756 54368 1820 54372
rect 99668 54428 99732 54432
rect 99668 54372 99672 54428
rect 99672 54372 99728 54428
rect 99728 54372 99732 54428
rect 99668 54368 99732 54372
rect 99748 54428 99812 54432
rect 99748 54372 99752 54428
rect 99752 54372 99808 54428
rect 99808 54372 99812 54428
rect 99748 54368 99812 54372
rect 99828 54428 99892 54432
rect 99828 54372 99832 54428
rect 99832 54372 99888 54428
rect 99888 54372 99892 54428
rect 99828 54368 99892 54372
rect 99908 54428 99972 54432
rect 99908 54372 99912 54428
rect 99912 54372 99968 54428
rect 99968 54372 99972 54428
rect 99908 54368 99972 54372
rect 1308 53884 1372 53888
rect 1308 53828 1312 53884
rect 1312 53828 1368 53884
rect 1368 53828 1372 53884
rect 1308 53824 1372 53828
rect 1388 53884 1452 53888
rect 1388 53828 1392 53884
rect 1392 53828 1448 53884
rect 1448 53828 1452 53884
rect 1388 53824 1452 53828
rect 98932 53884 98996 53888
rect 98932 53828 98936 53884
rect 98936 53828 98992 53884
rect 98992 53828 98996 53884
rect 98932 53824 98996 53828
rect 99012 53884 99076 53888
rect 99012 53828 99016 53884
rect 99016 53828 99072 53884
rect 99072 53828 99076 53884
rect 99012 53824 99076 53828
rect 99092 53884 99156 53888
rect 99092 53828 99096 53884
rect 99096 53828 99152 53884
rect 99152 53828 99156 53884
rect 99092 53824 99156 53828
rect 99172 53884 99236 53888
rect 99172 53828 99176 53884
rect 99176 53828 99232 53884
rect 99232 53828 99236 53884
rect 99172 53824 99236 53828
rect 1676 53340 1740 53344
rect 1676 53284 1680 53340
rect 1680 53284 1736 53340
rect 1736 53284 1740 53340
rect 1676 53280 1740 53284
rect 1756 53340 1820 53344
rect 1756 53284 1760 53340
rect 1760 53284 1816 53340
rect 1816 53284 1820 53340
rect 1756 53280 1820 53284
rect 99668 53340 99732 53344
rect 99668 53284 99672 53340
rect 99672 53284 99728 53340
rect 99728 53284 99732 53340
rect 99668 53280 99732 53284
rect 99748 53340 99812 53344
rect 99748 53284 99752 53340
rect 99752 53284 99808 53340
rect 99808 53284 99812 53340
rect 99748 53280 99812 53284
rect 99828 53340 99892 53344
rect 99828 53284 99832 53340
rect 99832 53284 99888 53340
rect 99888 53284 99892 53340
rect 99828 53280 99892 53284
rect 99908 53340 99972 53344
rect 99908 53284 99912 53340
rect 99912 53284 99968 53340
rect 99968 53284 99972 53340
rect 99908 53280 99972 53284
rect 1308 52796 1372 52800
rect 1308 52740 1312 52796
rect 1312 52740 1368 52796
rect 1368 52740 1372 52796
rect 1308 52736 1372 52740
rect 1388 52796 1452 52800
rect 1388 52740 1392 52796
rect 1392 52740 1448 52796
rect 1448 52740 1452 52796
rect 1388 52736 1452 52740
rect 98932 52796 98996 52800
rect 98932 52740 98936 52796
rect 98936 52740 98992 52796
rect 98992 52740 98996 52796
rect 98932 52736 98996 52740
rect 99012 52796 99076 52800
rect 99012 52740 99016 52796
rect 99016 52740 99072 52796
rect 99072 52740 99076 52796
rect 99012 52736 99076 52740
rect 99092 52796 99156 52800
rect 99092 52740 99096 52796
rect 99096 52740 99152 52796
rect 99152 52740 99156 52796
rect 99092 52736 99156 52740
rect 99172 52796 99236 52800
rect 99172 52740 99176 52796
rect 99176 52740 99232 52796
rect 99232 52740 99236 52796
rect 99172 52736 99236 52740
rect 1676 52252 1740 52256
rect 1676 52196 1680 52252
rect 1680 52196 1736 52252
rect 1736 52196 1740 52252
rect 1676 52192 1740 52196
rect 1756 52252 1820 52256
rect 1756 52196 1760 52252
rect 1760 52196 1816 52252
rect 1816 52196 1820 52252
rect 1756 52192 1820 52196
rect 99668 52252 99732 52256
rect 99668 52196 99672 52252
rect 99672 52196 99728 52252
rect 99728 52196 99732 52252
rect 99668 52192 99732 52196
rect 99748 52252 99812 52256
rect 99748 52196 99752 52252
rect 99752 52196 99808 52252
rect 99808 52196 99812 52252
rect 99748 52192 99812 52196
rect 99828 52252 99892 52256
rect 99828 52196 99832 52252
rect 99832 52196 99888 52252
rect 99888 52196 99892 52252
rect 99828 52192 99892 52196
rect 99908 52252 99972 52256
rect 99908 52196 99912 52252
rect 99912 52196 99968 52252
rect 99968 52196 99972 52252
rect 99908 52192 99972 52196
rect 1308 51708 1372 51712
rect 1308 51652 1312 51708
rect 1312 51652 1368 51708
rect 1368 51652 1372 51708
rect 1308 51648 1372 51652
rect 1388 51708 1452 51712
rect 1388 51652 1392 51708
rect 1392 51652 1448 51708
rect 1448 51652 1452 51708
rect 1388 51648 1452 51652
rect 98932 51708 98996 51712
rect 98932 51652 98936 51708
rect 98936 51652 98992 51708
rect 98992 51652 98996 51708
rect 98932 51648 98996 51652
rect 99012 51708 99076 51712
rect 99012 51652 99016 51708
rect 99016 51652 99072 51708
rect 99072 51652 99076 51708
rect 99012 51648 99076 51652
rect 99092 51708 99156 51712
rect 99092 51652 99096 51708
rect 99096 51652 99152 51708
rect 99152 51652 99156 51708
rect 99092 51648 99156 51652
rect 99172 51708 99236 51712
rect 99172 51652 99176 51708
rect 99176 51652 99232 51708
rect 99232 51652 99236 51708
rect 99172 51648 99236 51652
rect 1676 51164 1740 51168
rect 1676 51108 1680 51164
rect 1680 51108 1736 51164
rect 1736 51108 1740 51164
rect 1676 51104 1740 51108
rect 1756 51164 1820 51168
rect 1756 51108 1760 51164
rect 1760 51108 1816 51164
rect 1816 51108 1820 51164
rect 1756 51104 1820 51108
rect 99668 51164 99732 51168
rect 99668 51108 99672 51164
rect 99672 51108 99728 51164
rect 99728 51108 99732 51164
rect 99668 51104 99732 51108
rect 99748 51164 99812 51168
rect 99748 51108 99752 51164
rect 99752 51108 99808 51164
rect 99808 51108 99812 51164
rect 99748 51104 99812 51108
rect 99828 51164 99892 51168
rect 99828 51108 99832 51164
rect 99832 51108 99888 51164
rect 99888 51108 99892 51164
rect 99828 51104 99892 51108
rect 99908 51164 99972 51168
rect 99908 51108 99912 51164
rect 99912 51108 99968 51164
rect 99968 51108 99972 51164
rect 99908 51104 99972 51108
rect 1308 50620 1372 50624
rect 1308 50564 1312 50620
rect 1312 50564 1368 50620
rect 1368 50564 1372 50620
rect 1308 50560 1372 50564
rect 1388 50620 1452 50624
rect 1388 50564 1392 50620
rect 1392 50564 1448 50620
rect 1448 50564 1452 50620
rect 1388 50560 1452 50564
rect 98932 50620 98996 50624
rect 98932 50564 98936 50620
rect 98936 50564 98992 50620
rect 98992 50564 98996 50620
rect 98932 50560 98996 50564
rect 99012 50620 99076 50624
rect 99012 50564 99016 50620
rect 99016 50564 99072 50620
rect 99072 50564 99076 50620
rect 99012 50560 99076 50564
rect 99092 50620 99156 50624
rect 99092 50564 99096 50620
rect 99096 50564 99152 50620
rect 99152 50564 99156 50620
rect 99092 50560 99156 50564
rect 99172 50620 99236 50624
rect 99172 50564 99176 50620
rect 99176 50564 99232 50620
rect 99232 50564 99236 50620
rect 99172 50560 99236 50564
rect 1676 50076 1740 50080
rect 1676 50020 1680 50076
rect 1680 50020 1736 50076
rect 1736 50020 1740 50076
rect 1676 50016 1740 50020
rect 1756 50076 1820 50080
rect 1756 50020 1760 50076
rect 1760 50020 1816 50076
rect 1816 50020 1820 50076
rect 1756 50016 1820 50020
rect 99668 50076 99732 50080
rect 99668 50020 99672 50076
rect 99672 50020 99728 50076
rect 99728 50020 99732 50076
rect 99668 50016 99732 50020
rect 99748 50076 99812 50080
rect 99748 50020 99752 50076
rect 99752 50020 99808 50076
rect 99808 50020 99812 50076
rect 99748 50016 99812 50020
rect 99828 50076 99892 50080
rect 99828 50020 99832 50076
rect 99832 50020 99888 50076
rect 99888 50020 99892 50076
rect 99828 50016 99892 50020
rect 99908 50076 99972 50080
rect 99908 50020 99912 50076
rect 99912 50020 99968 50076
rect 99968 50020 99972 50076
rect 99908 50016 99972 50020
rect 1308 49532 1372 49536
rect 1308 49476 1312 49532
rect 1312 49476 1368 49532
rect 1368 49476 1372 49532
rect 1308 49472 1372 49476
rect 1388 49532 1452 49536
rect 1388 49476 1392 49532
rect 1392 49476 1448 49532
rect 1448 49476 1452 49532
rect 1388 49472 1452 49476
rect 98932 49532 98996 49536
rect 98932 49476 98936 49532
rect 98936 49476 98992 49532
rect 98992 49476 98996 49532
rect 98932 49472 98996 49476
rect 99012 49532 99076 49536
rect 99012 49476 99016 49532
rect 99016 49476 99072 49532
rect 99072 49476 99076 49532
rect 99012 49472 99076 49476
rect 99092 49532 99156 49536
rect 99092 49476 99096 49532
rect 99096 49476 99152 49532
rect 99152 49476 99156 49532
rect 99092 49472 99156 49476
rect 99172 49532 99236 49536
rect 99172 49476 99176 49532
rect 99176 49476 99232 49532
rect 99232 49476 99236 49532
rect 99172 49472 99236 49476
rect 1676 48988 1740 48992
rect 1676 48932 1680 48988
rect 1680 48932 1736 48988
rect 1736 48932 1740 48988
rect 1676 48928 1740 48932
rect 1756 48988 1820 48992
rect 1756 48932 1760 48988
rect 1760 48932 1816 48988
rect 1816 48932 1820 48988
rect 1756 48928 1820 48932
rect 99668 48988 99732 48992
rect 99668 48932 99672 48988
rect 99672 48932 99728 48988
rect 99728 48932 99732 48988
rect 99668 48928 99732 48932
rect 99748 48988 99812 48992
rect 99748 48932 99752 48988
rect 99752 48932 99808 48988
rect 99808 48932 99812 48988
rect 99748 48928 99812 48932
rect 99828 48988 99892 48992
rect 99828 48932 99832 48988
rect 99832 48932 99888 48988
rect 99888 48932 99892 48988
rect 99828 48928 99892 48932
rect 99908 48988 99972 48992
rect 99908 48932 99912 48988
rect 99912 48932 99968 48988
rect 99968 48932 99972 48988
rect 99908 48928 99972 48932
rect 1308 48444 1372 48448
rect 1308 48388 1312 48444
rect 1312 48388 1368 48444
rect 1368 48388 1372 48444
rect 1308 48384 1372 48388
rect 1388 48444 1452 48448
rect 1388 48388 1392 48444
rect 1392 48388 1448 48444
rect 1448 48388 1452 48444
rect 1388 48384 1452 48388
rect 98932 48444 98996 48448
rect 98932 48388 98936 48444
rect 98936 48388 98992 48444
rect 98992 48388 98996 48444
rect 98932 48384 98996 48388
rect 99012 48444 99076 48448
rect 99012 48388 99016 48444
rect 99016 48388 99072 48444
rect 99072 48388 99076 48444
rect 99012 48384 99076 48388
rect 99092 48444 99156 48448
rect 99092 48388 99096 48444
rect 99096 48388 99152 48444
rect 99152 48388 99156 48444
rect 99092 48384 99156 48388
rect 99172 48444 99236 48448
rect 99172 48388 99176 48444
rect 99176 48388 99232 48444
rect 99232 48388 99236 48444
rect 99172 48384 99236 48388
rect 1676 47900 1740 47904
rect 1676 47844 1680 47900
rect 1680 47844 1736 47900
rect 1736 47844 1740 47900
rect 1676 47840 1740 47844
rect 1756 47900 1820 47904
rect 1756 47844 1760 47900
rect 1760 47844 1816 47900
rect 1816 47844 1820 47900
rect 1756 47840 1820 47844
rect 99668 47900 99732 47904
rect 99668 47844 99672 47900
rect 99672 47844 99728 47900
rect 99728 47844 99732 47900
rect 99668 47840 99732 47844
rect 99748 47900 99812 47904
rect 99748 47844 99752 47900
rect 99752 47844 99808 47900
rect 99808 47844 99812 47900
rect 99748 47840 99812 47844
rect 99828 47900 99892 47904
rect 99828 47844 99832 47900
rect 99832 47844 99888 47900
rect 99888 47844 99892 47900
rect 99828 47840 99892 47844
rect 99908 47900 99972 47904
rect 99908 47844 99912 47900
rect 99912 47844 99968 47900
rect 99968 47844 99972 47900
rect 99908 47840 99972 47844
rect 1308 47356 1372 47360
rect 1308 47300 1312 47356
rect 1312 47300 1368 47356
rect 1368 47300 1372 47356
rect 1308 47296 1372 47300
rect 1388 47356 1452 47360
rect 1388 47300 1392 47356
rect 1392 47300 1448 47356
rect 1448 47300 1452 47356
rect 1388 47296 1452 47300
rect 98932 47356 98996 47360
rect 98932 47300 98936 47356
rect 98936 47300 98992 47356
rect 98992 47300 98996 47356
rect 98932 47296 98996 47300
rect 99012 47356 99076 47360
rect 99012 47300 99016 47356
rect 99016 47300 99072 47356
rect 99072 47300 99076 47356
rect 99012 47296 99076 47300
rect 99092 47356 99156 47360
rect 99092 47300 99096 47356
rect 99096 47300 99152 47356
rect 99152 47300 99156 47356
rect 99092 47296 99156 47300
rect 99172 47356 99236 47360
rect 99172 47300 99176 47356
rect 99176 47300 99232 47356
rect 99232 47300 99236 47356
rect 99172 47296 99236 47300
rect 1676 46812 1740 46816
rect 1676 46756 1680 46812
rect 1680 46756 1736 46812
rect 1736 46756 1740 46812
rect 1676 46752 1740 46756
rect 1756 46812 1820 46816
rect 1756 46756 1760 46812
rect 1760 46756 1816 46812
rect 1816 46756 1820 46812
rect 1756 46752 1820 46756
rect 99668 46812 99732 46816
rect 99668 46756 99672 46812
rect 99672 46756 99728 46812
rect 99728 46756 99732 46812
rect 99668 46752 99732 46756
rect 99748 46812 99812 46816
rect 99748 46756 99752 46812
rect 99752 46756 99808 46812
rect 99808 46756 99812 46812
rect 99748 46752 99812 46756
rect 99828 46812 99892 46816
rect 99828 46756 99832 46812
rect 99832 46756 99888 46812
rect 99888 46756 99892 46812
rect 99828 46752 99892 46756
rect 99908 46812 99972 46816
rect 99908 46756 99912 46812
rect 99912 46756 99968 46812
rect 99968 46756 99972 46812
rect 99908 46752 99972 46756
rect 1308 46268 1372 46272
rect 1308 46212 1312 46268
rect 1312 46212 1368 46268
rect 1368 46212 1372 46268
rect 1308 46208 1372 46212
rect 1388 46268 1452 46272
rect 1388 46212 1392 46268
rect 1392 46212 1448 46268
rect 1448 46212 1452 46268
rect 1388 46208 1452 46212
rect 98932 46268 98996 46272
rect 98932 46212 98936 46268
rect 98936 46212 98992 46268
rect 98992 46212 98996 46268
rect 98932 46208 98996 46212
rect 99012 46268 99076 46272
rect 99012 46212 99016 46268
rect 99016 46212 99072 46268
rect 99072 46212 99076 46268
rect 99012 46208 99076 46212
rect 99092 46268 99156 46272
rect 99092 46212 99096 46268
rect 99096 46212 99152 46268
rect 99152 46212 99156 46268
rect 99092 46208 99156 46212
rect 99172 46268 99236 46272
rect 99172 46212 99176 46268
rect 99176 46212 99232 46268
rect 99232 46212 99236 46268
rect 99172 46208 99236 46212
rect 1676 45724 1740 45728
rect 1676 45668 1680 45724
rect 1680 45668 1736 45724
rect 1736 45668 1740 45724
rect 1676 45664 1740 45668
rect 1756 45724 1820 45728
rect 1756 45668 1760 45724
rect 1760 45668 1816 45724
rect 1816 45668 1820 45724
rect 1756 45664 1820 45668
rect 99668 45724 99732 45728
rect 99668 45668 99672 45724
rect 99672 45668 99728 45724
rect 99728 45668 99732 45724
rect 99668 45664 99732 45668
rect 99748 45724 99812 45728
rect 99748 45668 99752 45724
rect 99752 45668 99808 45724
rect 99808 45668 99812 45724
rect 99748 45664 99812 45668
rect 99828 45724 99892 45728
rect 99828 45668 99832 45724
rect 99832 45668 99888 45724
rect 99888 45668 99892 45724
rect 99828 45664 99892 45668
rect 99908 45724 99972 45728
rect 99908 45668 99912 45724
rect 99912 45668 99968 45724
rect 99968 45668 99972 45724
rect 99908 45664 99972 45668
rect 1308 45180 1372 45184
rect 1308 45124 1312 45180
rect 1312 45124 1368 45180
rect 1368 45124 1372 45180
rect 1308 45120 1372 45124
rect 1388 45180 1452 45184
rect 1388 45124 1392 45180
rect 1392 45124 1448 45180
rect 1448 45124 1452 45180
rect 1388 45120 1452 45124
rect 98932 45180 98996 45184
rect 98932 45124 98936 45180
rect 98936 45124 98992 45180
rect 98992 45124 98996 45180
rect 98932 45120 98996 45124
rect 99012 45180 99076 45184
rect 99012 45124 99016 45180
rect 99016 45124 99072 45180
rect 99072 45124 99076 45180
rect 99012 45120 99076 45124
rect 99092 45180 99156 45184
rect 99092 45124 99096 45180
rect 99096 45124 99152 45180
rect 99152 45124 99156 45180
rect 99092 45120 99156 45124
rect 99172 45180 99236 45184
rect 99172 45124 99176 45180
rect 99176 45124 99232 45180
rect 99232 45124 99236 45180
rect 99172 45120 99236 45124
rect 1676 44636 1740 44640
rect 1676 44580 1680 44636
rect 1680 44580 1736 44636
rect 1736 44580 1740 44636
rect 1676 44576 1740 44580
rect 1756 44636 1820 44640
rect 1756 44580 1760 44636
rect 1760 44580 1816 44636
rect 1816 44580 1820 44636
rect 1756 44576 1820 44580
rect 99668 44636 99732 44640
rect 99668 44580 99672 44636
rect 99672 44580 99728 44636
rect 99728 44580 99732 44636
rect 99668 44576 99732 44580
rect 99748 44636 99812 44640
rect 99748 44580 99752 44636
rect 99752 44580 99808 44636
rect 99808 44580 99812 44636
rect 99748 44576 99812 44580
rect 99828 44636 99892 44640
rect 99828 44580 99832 44636
rect 99832 44580 99888 44636
rect 99888 44580 99892 44636
rect 99828 44576 99892 44580
rect 99908 44636 99972 44640
rect 99908 44580 99912 44636
rect 99912 44580 99968 44636
rect 99968 44580 99972 44636
rect 99908 44576 99972 44580
rect 1308 44092 1372 44096
rect 1308 44036 1312 44092
rect 1312 44036 1368 44092
rect 1368 44036 1372 44092
rect 1308 44032 1372 44036
rect 1388 44092 1452 44096
rect 1388 44036 1392 44092
rect 1392 44036 1448 44092
rect 1448 44036 1452 44092
rect 1388 44032 1452 44036
rect 98932 44092 98996 44096
rect 98932 44036 98936 44092
rect 98936 44036 98992 44092
rect 98992 44036 98996 44092
rect 98932 44032 98996 44036
rect 99012 44092 99076 44096
rect 99012 44036 99016 44092
rect 99016 44036 99072 44092
rect 99072 44036 99076 44092
rect 99012 44032 99076 44036
rect 99092 44092 99156 44096
rect 99092 44036 99096 44092
rect 99096 44036 99152 44092
rect 99152 44036 99156 44092
rect 99092 44032 99156 44036
rect 99172 44092 99236 44096
rect 99172 44036 99176 44092
rect 99176 44036 99232 44092
rect 99232 44036 99236 44092
rect 99172 44032 99236 44036
rect 1676 43548 1740 43552
rect 1676 43492 1680 43548
rect 1680 43492 1736 43548
rect 1736 43492 1740 43548
rect 1676 43488 1740 43492
rect 1756 43548 1820 43552
rect 1756 43492 1760 43548
rect 1760 43492 1816 43548
rect 1816 43492 1820 43548
rect 1756 43488 1820 43492
rect 99668 43548 99732 43552
rect 99668 43492 99672 43548
rect 99672 43492 99728 43548
rect 99728 43492 99732 43548
rect 99668 43488 99732 43492
rect 99748 43548 99812 43552
rect 99748 43492 99752 43548
rect 99752 43492 99808 43548
rect 99808 43492 99812 43548
rect 99748 43488 99812 43492
rect 99828 43548 99892 43552
rect 99828 43492 99832 43548
rect 99832 43492 99888 43548
rect 99888 43492 99892 43548
rect 99828 43488 99892 43492
rect 99908 43548 99972 43552
rect 99908 43492 99912 43548
rect 99912 43492 99968 43548
rect 99968 43492 99972 43548
rect 99908 43488 99972 43492
rect 1308 43004 1372 43008
rect 1308 42948 1312 43004
rect 1312 42948 1368 43004
rect 1368 42948 1372 43004
rect 1308 42944 1372 42948
rect 1388 43004 1452 43008
rect 1388 42948 1392 43004
rect 1392 42948 1448 43004
rect 1448 42948 1452 43004
rect 1388 42944 1452 42948
rect 98932 43004 98996 43008
rect 98932 42948 98936 43004
rect 98936 42948 98992 43004
rect 98992 42948 98996 43004
rect 98932 42944 98996 42948
rect 99012 43004 99076 43008
rect 99012 42948 99016 43004
rect 99016 42948 99072 43004
rect 99072 42948 99076 43004
rect 99012 42944 99076 42948
rect 99092 43004 99156 43008
rect 99092 42948 99096 43004
rect 99096 42948 99152 43004
rect 99152 42948 99156 43004
rect 99092 42944 99156 42948
rect 99172 43004 99236 43008
rect 99172 42948 99176 43004
rect 99176 42948 99232 43004
rect 99232 42948 99236 43004
rect 99172 42944 99236 42948
rect 1676 42460 1740 42464
rect 1676 42404 1680 42460
rect 1680 42404 1736 42460
rect 1736 42404 1740 42460
rect 1676 42400 1740 42404
rect 1756 42460 1820 42464
rect 1756 42404 1760 42460
rect 1760 42404 1816 42460
rect 1816 42404 1820 42460
rect 1756 42400 1820 42404
rect 99668 42460 99732 42464
rect 99668 42404 99672 42460
rect 99672 42404 99728 42460
rect 99728 42404 99732 42460
rect 99668 42400 99732 42404
rect 99748 42460 99812 42464
rect 99748 42404 99752 42460
rect 99752 42404 99808 42460
rect 99808 42404 99812 42460
rect 99748 42400 99812 42404
rect 99828 42460 99892 42464
rect 99828 42404 99832 42460
rect 99832 42404 99888 42460
rect 99888 42404 99892 42460
rect 99828 42400 99892 42404
rect 99908 42460 99972 42464
rect 99908 42404 99912 42460
rect 99912 42404 99968 42460
rect 99968 42404 99972 42460
rect 99908 42400 99972 42404
rect 1308 41916 1372 41920
rect 1308 41860 1312 41916
rect 1312 41860 1368 41916
rect 1368 41860 1372 41916
rect 1308 41856 1372 41860
rect 1388 41916 1452 41920
rect 1388 41860 1392 41916
rect 1392 41860 1448 41916
rect 1448 41860 1452 41916
rect 1388 41856 1452 41860
rect 98932 41916 98996 41920
rect 98932 41860 98936 41916
rect 98936 41860 98992 41916
rect 98992 41860 98996 41916
rect 98932 41856 98996 41860
rect 99012 41916 99076 41920
rect 99012 41860 99016 41916
rect 99016 41860 99072 41916
rect 99072 41860 99076 41916
rect 99012 41856 99076 41860
rect 99092 41916 99156 41920
rect 99092 41860 99096 41916
rect 99096 41860 99152 41916
rect 99152 41860 99156 41916
rect 99092 41856 99156 41860
rect 99172 41916 99236 41920
rect 99172 41860 99176 41916
rect 99176 41860 99232 41916
rect 99232 41860 99236 41916
rect 99172 41856 99236 41860
rect 1676 41372 1740 41376
rect 1676 41316 1680 41372
rect 1680 41316 1736 41372
rect 1736 41316 1740 41372
rect 1676 41312 1740 41316
rect 1756 41372 1820 41376
rect 1756 41316 1760 41372
rect 1760 41316 1816 41372
rect 1816 41316 1820 41372
rect 1756 41312 1820 41316
rect 99668 41372 99732 41376
rect 99668 41316 99672 41372
rect 99672 41316 99728 41372
rect 99728 41316 99732 41372
rect 99668 41312 99732 41316
rect 99748 41372 99812 41376
rect 99748 41316 99752 41372
rect 99752 41316 99808 41372
rect 99808 41316 99812 41372
rect 99748 41312 99812 41316
rect 99828 41372 99892 41376
rect 99828 41316 99832 41372
rect 99832 41316 99888 41372
rect 99888 41316 99892 41372
rect 99828 41312 99892 41316
rect 99908 41372 99972 41376
rect 99908 41316 99912 41372
rect 99912 41316 99968 41372
rect 99968 41316 99972 41372
rect 99908 41312 99972 41316
rect 1308 40828 1372 40832
rect 1308 40772 1312 40828
rect 1312 40772 1368 40828
rect 1368 40772 1372 40828
rect 1308 40768 1372 40772
rect 1388 40828 1452 40832
rect 1388 40772 1392 40828
rect 1392 40772 1448 40828
rect 1448 40772 1452 40828
rect 1388 40768 1452 40772
rect 98932 40828 98996 40832
rect 98932 40772 98936 40828
rect 98936 40772 98992 40828
rect 98992 40772 98996 40828
rect 98932 40768 98996 40772
rect 99012 40828 99076 40832
rect 99012 40772 99016 40828
rect 99016 40772 99072 40828
rect 99072 40772 99076 40828
rect 99012 40768 99076 40772
rect 99092 40828 99156 40832
rect 99092 40772 99096 40828
rect 99096 40772 99152 40828
rect 99152 40772 99156 40828
rect 99092 40768 99156 40772
rect 99172 40828 99236 40832
rect 99172 40772 99176 40828
rect 99176 40772 99232 40828
rect 99232 40772 99236 40828
rect 99172 40768 99236 40772
rect 1676 40284 1740 40288
rect 1676 40228 1680 40284
rect 1680 40228 1736 40284
rect 1736 40228 1740 40284
rect 1676 40224 1740 40228
rect 1756 40284 1820 40288
rect 1756 40228 1760 40284
rect 1760 40228 1816 40284
rect 1816 40228 1820 40284
rect 1756 40224 1820 40228
rect 99668 40284 99732 40288
rect 99668 40228 99672 40284
rect 99672 40228 99728 40284
rect 99728 40228 99732 40284
rect 99668 40224 99732 40228
rect 99748 40284 99812 40288
rect 99748 40228 99752 40284
rect 99752 40228 99808 40284
rect 99808 40228 99812 40284
rect 99748 40224 99812 40228
rect 99828 40284 99892 40288
rect 99828 40228 99832 40284
rect 99832 40228 99888 40284
rect 99888 40228 99892 40284
rect 99828 40224 99892 40228
rect 99908 40284 99972 40288
rect 99908 40228 99912 40284
rect 99912 40228 99968 40284
rect 99968 40228 99972 40284
rect 99908 40224 99972 40228
rect 1308 39740 1372 39744
rect 1308 39684 1312 39740
rect 1312 39684 1368 39740
rect 1368 39684 1372 39740
rect 1308 39680 1372 39684
rect 1388 39740 1452 39744
rect 1388 39684 1392 39740
rect 1392 39684 1448 39740
rect 1448 39684 1452 39740
rect 1388 39680 1452 39684
rect 98932 39740 98996 39744
rect 98932 39684 98936 39740
rect 98936 39684 98992 39740
rect 98992 39684 98996 39740
rect 98932 39680 98996 39684
rect 99012 39740 99076 39744
rect 99012 39684 99016 39740
rect 99016 39684 99072 39740
rect 99072 39684 99076 39740
rect 99012 39680 99076 39684
rect 99092 39740 99156 39744
rect 99092 39684 99096 39740
rect 99096 39684 99152 39740
rect 99152 39684 99156 39740
rect 99092 39680 99156 39684
rect 99172 39740 99236 39744
rect 99172 39684 99176 39740
rect 99176 39684 99232 39740
rect 99232 39684 99236 39740
rect 99172 39680 99236 39684
rect 1676 39196 1740 39200
rect 1676 39140 1680 39196
rect 1680 39140 1736 39196
rect 1736 39140 1740 39196
rect 1676 39136 1740 39140
rect 1756 39196 1820 39200
rect 1756 39140 1760 39196
rect 1760 39140 1816 39196
rect 1816 39140 1820 39196
rect 1756 39136 1820 39140
rect 99668 39196 99732 39200
rect 99668 39140 99672 39196
rect 99672 39140 99728 39196
rect 99728 39140 99732 39196
rect 99668 39136 99732 39140
rect 99748 39196 99812 39200
rect 99748 39140 99752 39196
rect 99752 39140 99808 39196
rect 99808 39140 99812 39196
rect 99748 39136 99812 39140
rect 99828 39196 99892 39200
rect 99828 39140 99832 39196
rect 99832 39140 99888 39196
rect 99888 39140 99892 39196
rect 99828 39136 99892 39140
rect 99908 39196 99972 39200
rect 99908 39140 99912 39196
rect 99912 39140 99968 39196
rect 99968 39140 99972 39196
rect 99908 39136 99972 39140
rect 1308 38652 1372 38656
rect 1308 38596 1312 38652
rect 1312 38596 1368 38652
rect 1368 38596 1372 38652
rect 1308 38592 1372 38596
rect 1388 38652 1452 38656
rect 1388 38596 1392 38652
rect 1392 38596 1448 38652
rect 1448 38596 1452 38652
rect 1388 38592 1452 38596
rect 98932 38652 98996 38656
rect 98932 38596 98936 38652
rect 98936 38596 98992 38652
rect 98992 38596 98996 38652
rect 98932 38592 98996 38596
rect 99012 38652 99076 38656
rect 99012 38596 99016 38652
rect 99016 38596 99072 38652
rect 99072 38596 99076 38652
rect 99012 38592 99076 38596
rect 99092 38652 99156 38656
rect 99092 38596 99096 38652
rect 99096 38596 99152 38652
rect 99152 38596 99156 38652
rect 99092 38592 99156 38596
rect 99172 38652 99236 38656
rect 99172 38596 99176 38652
rect 99176 38596 99232 38652
rect 99232 38596 99236 38652
rect 99172 38592 99236 38596
rect 1676 38108 1740 38112
rect 1676 38052 1680 38108
rect 1680 38052 1736 38108
rect 1736 38052 1740 38108
rect 1676 38048 1740 38052
rect 1756 38108 1820 38112
rect 1756 38052 1760 38108
rect 1760 38052 1816 38108
rect 1816 38052 1820 38108
rect 1756 38048 1820 38052
rect 99668 38108 99732 38112
rect 99668 38052 99672 38108
rect 99672 38052 99728 38108
rect 99728 38052 99732 38108
rect 99668 38048 99732 38052
rect 99748 38108 99812 38112
rect 99748 38052 99752 38108
rect 99752 38052 99808 38108
rect 99808 38052 99812 38108
rect 99748 38048 99812 38052
rect 99828 38108 99892 38112
rect 99828 38052 99832 38108
rect 99832 38052 99888 38108
rect 99888 38052 99892 38108
rect 99828 38048 99892 38052
rect 99908 38108 99972 38112
rect 99908 38052 99912 38108
rect 99912 38052 99968 38108
rect 99968 38052 99972 38108
rect 99908 38048 99972 38052
rect 1308 37564 1372 37568
rect 1308 37508 1312 37564
rect 1312 37508 1368 37564
rect 1368 37508 1372 37564
rect 1308 37504 1372 37508
rect 1388 37564 1452 37568
rect 1388 37508 1392 37564
rect 1392 37508 1448 37564
rect 1448 37508 1452 37564
rect 1388 37504 1452 37508
rect 98932 37564 98996 37568
rect 98932 37508 98936 37564
rect 98936 37508 98992 37564
rect 98992 37508 98996 37564
rect 98932 37504 98996 37508
rect 99012 37564 99076 37568
rect 99012 37508 99016 37564
rect 99016 37508 99072 37564
rect 99072 37508 99076 37564
rect 99012 37504 99076 37508
rect 99092 37564 99156 37568
rect 99092 37508 99096 37564
rect 99096 37508 99152 37564
rect 99152 37508 99156 37564
rect 99092 37504 99156 37508
rect 99172 37564 99236 37568
rect 99172 37508 99176 37564
rect 99176 37508 99232 37564
rect 99232 37508 99236 37564
rect 99172 37504 99236 37508
rect 1676 37020 1740 37024
rect 1676 36964 1680 37020
rect 1680 36964 1736 37020
rect 1736 36964 1740 37020
rect 1676 36960 1740 36964
rect 1756 37020 1820 37024
rect 1756 36964 1760 37020
rect 1760 36964 1816 37020
rect 1816 36964 1820 37020
rect 1756 36960 1820 36964
rect 99668 37020 99732 37024
rect 99668 36964 99672 37020
rect 99672 36964 99728 37020
rect 99728 36964 99732 37020
rect 99668 36960 99732 36964
rect 99748 37020 99812 37024
rect 99748 36964 99752 37020
rect 99752 36964 99808 37020
rect 99808 36964 99812 37020
rect 99748 36960 99812 36964
rect 99828 37020 99892 37024
rect 99828 36964 99832 37020
rect 99832 36964 99888 37020
rect 99888 36964 99892 37020
rect 99828 36960 99892 36964
rect 99908 37020 99972 37024
rect 99908 36964 99912 37020
rect 99912 36964 99968 37020
rect 99968 36964 99972 37020
rect 99908 36960 99972 36964
rect 1308 36476 1372 36480
rect 1308 36420 1312 36476
rect 1312 36420 1368 36476
rect 1368 36420 1372 36476
rect 1308 36416 1372 36420
rect 1388 36476 1452 36480
rect 1388 36420 1392 36476
rect 1392 36420 1448 36476
rect 1448 36420 1452 36476
rect 1388 36416 1452 36420
rect 98932 36476 98996 36480
rect 98932 36420 98936 36476
rect 98936 36420 98992 36476
rect 98992 36420 98996 36476
rect 98932 36416 98996 36420
rect 99012 36476 99076 36480
rect 99012 36420 99016 36476
rect 99016 36420 99072 36476
rect 99072 36420 99076 36476
rect 99012 36416 99076 36420
rect 99092 36476 99156 36480
rect 99092 36420 99096 36476
rect 99096 36420 99152 36476
rect 99152 36420 99156 36476
rect 99092 36416 99156 36420
rect 99172 36476 99236 36480
rect 99172 36420 99176 36476
rect 99176 36420 99232 36476
rect 99232 36420 99236 36476
rect 99172 36416 99236 36420
rect 1676 35932 1740 35936
rect 1676 35876 1680 35932
rect 1680 35876 1736 35932
rect 1736 35876 1740 35932
rect 1676 35872 1740 35876
rect 1756 35932 1820 35936
rect 1756 35876 1760 35932
rect 1760 35876 1816 35932
rect 1816 35876 1820 35932
rect 1756 35872 1820 35876
rect 99668 35932 99732 35936
rect 99668 35876 99672 35932
rect 99672 35876 99728 35932
rect 99728 35876 99732 35932
rect 99668 35872 99732 35876
rect 99748 35932 99812 35936
rect 99748 35876 99752 35932
rect 99752 35876 99808 35932
rect 99808 35876 99812 35932
rect 99748 35872 99812 35876
rect 99828 35932 99892 35936
rect 99828 35876 99832 35932
rect 99832 35876 99888 35932
rect 99888 35876 99892 35932
rect 99828 35872 99892 35876
rect 99908 35932 99972 35936
rect 99908 35876 99912 35932
rect 99912 35876 99968 35932
rect 99968 35876 99972 35932
rect 99908 35872 99972 35876
rect 1308 35388 1372 35392
rect 1308 35332 1312 35388
rect 1312 35332 1368 35388
rect 1368 35332 1372 35388
rect 1308 35328 1372 35332
rect 1388 35388 1452 35392
rect 1388 35332 1392 35388
rect 1392 35332 1448 35388
rect 1448 35332 1452 35388
rect 1388 35328 1452 35332
rect 98932 35388 98996 35392
rect 98932 35332 98936 35388
rect 98936 35332 98992 35388
rect 98992 35332 98996 35388
rect 98932 35328 98996 35332
rect 99012 35388 99076 35392
rect 99012 35332 99016 35388
rect 99016 35332 99072 35388
rect 99072 35332 99076 35388
rect 99012 35328 99076 35332
rect 99092 35388 99156 35392
rect 99092 35332 99096 35388
rect 99096 35332 99152 35388
rect 99152 35332 99156 35388
rect 99092 35328 99156 35332
rect 99172 35388 99236 35392
rect 99172 35332 99176 35388
rect 99176 35332 99232 35388
rect 99232 35332 99236 35388
rect 99172 35328 99236 35332
rect 1676 34844 1740 34848
rect 1676 34788 1680 34844
rect 1680 34788 1736 34844
rect 1736 34788 1740 34844
rect 1676 34784 1740 34788
rect 1756 34844 1820 34848
rect 1756 34788 1760 34844
rect 1760 34788 1816 34844
rect 1816 34788 1820 34844
rect 1756 34784 1820 34788
rect 99668 34844 99732 34848
rect 99668 34788 99672 34844
rect 99672 34788 99728 34844
rect 99728 34788 99732 34844
rect 99668 34784 99732 34788
rect 99748 34844 99812 34848
rect 99748 34788 99752 34844
rect 99752 34788 99808 34844
rect 99808 34788 99812 34844
rect 99748 34784 99812 34788
rect 99828 34844 99892 34848
rect 99828 34788 99832 34844
rect 99832 34788 99888 34844
rect 99888 34788 99892 34844
rect 99828 34784 99892 34788
rect 99908 34844 99972 34848
rect 99908 34788 99912 34844
rect 99912 34788 99968 34844
rect 99968 34788 99972 34844
rect 99908 34784 99972 34788
rect 1308 34300 1372 34304
rect 1308 34244 1312 34300
rect 1312 34244 1368 34300
rect 1368 34244 1372 34300
rect 1308 34240 1372 34244
rect 1388 34300 1452 34304
rect 1388 34244 1392 34300
rect 1392 34244 1448 34300
rect 1448 34244 1452 34300
rect 1388 34240 1452 34244
rect 98932 34300 98996 34304
rect 98932 34244 98936 34300
rect 98936 34244 98992 34300
rect 98992 34244 98996 34300
rect 98932 34240 98996 34244
rect 99012 34300 99076 34304
rect 99012 34244 99016 34300
rect 99016 34244 99072 34300
rect 99072 34244 99076 34300
rect 99012 34240 99076 34244
rect 99092 34300 99156 34304
rect 99092 34244 99096 34300
rect 99096 34244 99152 34300
rect 99152 34244 99156 34300
rect 99092 34240 99156 34244
rect 99172 34300 99236 34304
rect 99172 34244 99176 34300
rect 99176 34244 99232 34300
rect 99232 34244 99236 34300
rect 99172 34240 99236 34244
rect 1676 33756 1740 33760
rect 1676 33700 1680 33756
rect 1680 33700 1736 33756
rect 1736 33700 1740 33756
rect 1676 33696 1740 33700
rect 1756 33756 1820 33760
rect 1756 33700 1760 33756
rect 1760 33700 1816 33756
rect 1816 33700 1820 33756
rect 1756 33696 1820 33700
rect 99668 33756 99732 33760
rect 99668 33700 99672 33756
rect 99672 33700 99728 33756
rect 99728 33700 99732 33756
rect 99668 33696 99732 33700
rect 99748 33756 99812 33760
rect 99748 33700 99752 33756
rect 99752 33700 99808 33756
rect 99808 33700 99812 33756
rect 99748 33696 99812 33700
rect 99828 33756 99892 33760
rect 99828 33700 99832 33756
rect 99832 33700 99888 33756
rect 99888 33700 99892 33756
rect 99828 33696 99892 33700
rect 99908 33756 99972 33760
rect 99908 33700 99912 33756
rect 99912 33700 99968 33756
rect 99968 33700 99972 33756
rect 99908 33696 99972 33700
rect 1308 33212 1372 33216
rect 1308 33156 1312 33212
rect 1312 33156 1368 33212
rect 1368 33156 1372 33212
rect 1308 33152 1372 33156
rect 1388 33212 1452 33216
rect 1388 33156 1392 33212
rect 1392 33156 1448 33212
rect 1448 33156 1452 33212
rect 1388 33152 1452 33156
rect 98932 33212 98996 33216
rect 98932 33156 98936 33212
rect 98936 33156 98992 33212
rect 98992 33156 98996 33212
rect 98932 33152 98996 33156
rect 99012 33212 99076 33216
rect 99012 33156 99016 33212
rect 99016 33156 99072 33212
rect 99072 33156 99076 33212
rect 99012 33152 99076 33156
rect 99092 33212 99156 33216
rect 99092 33156 99096 33212
rect 99096 33156 99152 33212
rect 99152 33156 99156 33212
rect 99092 33152 99156 33156
rect 99172 33212 99236 33216
rect 99172 33156 99176 33212
rect 99176 33156 99232 33212
rect 99232 33156 99236 33212
rect 99172 33152 99236 33156
rect 1676 32668 1740 32672
rect 1676 32612 1680 32668
rect 1680 32612 1736 32668
rect 1736 32612 1740 32668
rect 1676 32608 1740 32612
rect 1756 32668 1820 32672
rect 1756 32612 1760 32668
rect 1760 32612 1816 32668
rect 1816 32612 1820 32668
rect 1756 32608 1820 32612
rect 99668 32668 99732 32672
rect 99668 32612 99672 32668
rect 99672 32612 99728 32668
rect 99728 32612 99732 32668
rect 99668 32608 99732 32612
rect 99748 32668 99812 32672
rect 99748 32612 99752 32668
rect 99752 32612 99808 32668
rect 99808 32612 99812 32668
rect 99748 32608 99812 32612
rect 99828 32668 99892 32672
rect 99828 32612 99832 32668
rect 99832 32612 99888 32668
rect 99888 32612 99892 32668
rect 99828 32608 99892 32612
rect 99908 32668 99972 32672
rect 99908 32612 99912 32668
rect 99912 32612 99968 32668
rect 99968 32612 99972 32668
rect 99908 32608 99972 32612
rect 1308 32124 1372 32128
rect 1308 32068 1312 32124
rect 1312 32068 1368 32124
rect 1368 32068 1372 32124
rect 1308 32064 1372 32068
rect 1388 32124 1452 32128
rect 1388 32068 1392 32124
rect 1392 32068 1448 32124
rect 1448 32068 1452 32124
rect 1388 32064 1452 32068
rect 98932 32124 98996 32128
rect 98932 32068 98936 32124
rect 98936 32068 98992 32124
rect 98992 32068 98996 32124
rect 98932 32064 98996 32068
rect 99012 32124 99076 32128
rect 99012 32068 99016 32124
rect 99016 32068 99072 32124
rect 99072 32068 99076 32124
rect 99012 32064 99076 32068
rect 99092 32124 99156 32128
rect 99092 32068 99096 32124
rect 99096 32068 99152 32124
rect 99152 32068 99156 32124
rect 99092 32064 99156 32068
rect 99172 32124 99236 32128
rect 99172 32068 99176 32124
rect 99176 32068 99232 32124
rect 99232 32068 99236 32124
rect 99172 32064 99236 32068
rect 1676 31580 1740 31584
rect 1676 31524 1680 31580
rect 1680 31524 1736 31580
rect 1736 31524 1740 31580
rect 1676 31520 1740 31524
rect 1756 31580 1820 31584
rect 1756 31524 1760 31580
rect 1760 31524 1816 31580
rect 1816 31524 1820 31580
rect 1756 31520 1820 31524
rect 99668 31580 99732 31584
rect 99668 31524 99672 31580
rect 99672 31524 99728 31580
rect 99728 31524 99732 31580
rect 99668 31520 99732 31524
rect 99748 31580 99812 31584
rect 99748 31524 99752 31580
rect 99752 31524 99808 31580
rect 99808 31524 99812 31580
rect 99748 31520 99812 31524
rect 99828 31580 99892 31584
rect 99828 31524 99832 31580
rect 99832 31524 99888 31580
rect 99888 31524 99892 31580
rect 99828 31520 99892 31524
rect 99908 31580 99972 31584
rect 99908 31524 99912 31580
rect 99912 31524 99968 31580
rect 99968 31524 99972 31580
rect 99908 31520 99972 31524
rect 1308 31036 1372 31040
rect 1308 30980 1312 31036
rect 1312 30980 1368 31036
rect 1368 30980 1372 31036
rect 1308 30976 1372 30980
rect 1388 31036 1452 31040
rect 1388 30980 1392 31036
rect 1392 30980 1448 31036
rect 1448 30980 1452 31036
rect 1388 30976 1452 30980
rect 98932 31036 98996 31040
rect 98932 30980 98936 31036
rect 98936 30980 98992 31036
rect 98992 30980 98996 31036
rect 98932 30976 98996 30980
rect 99012 31036 99076 31040
rect 99012 30980 99016 31036
rect 99016 30980 99072 31036
rect 99072 30980 99076 31036
rect 99012 30976 99076 30980
rect 99092 31036 99156 31040
rect 99092 30980 99096 31036
rect 99096 30980 99152 31036
rect 99152 30980 99156 31036
rect 99092 30976 99156 30980
rect 99172 31036 99236 31040
rect 99172 30980 99176 31036
rect 99176 30980 99232 31036
rect 99232 30980 99236 31036
rect 99172 30976 99236 30980
rect 1676 30492 1740 30496
rect 1676 30436 1680 30492
rect 1680 30436 1736 30492
rect 1736 30436 1740 30492
rect 1676 30432 1740 30436
rect 1756 30492 1820 30496
rect 1756 30436 1760 30492
rect 1760 30436 1816 30492
rect 1816 30436 1820 30492
rect 1756 30432 1820 30436
rect 99668 30492 99732 30496
rect 99668 30436 99672 30492
rect 99672 30436 99728 30492
rect 99728 30436 99732 30492
rect 99668 30432 99732 30436
rect 99748 30492 99812 30496
rect 99748 30436 99752 30492
rect 99752 30436 99808 30492
rect 99808 30436 99812 30492
rect 99748 30432 99812 30436
rect 99828 30492 99892 30496
rect 99828 30436 99832 30492
rect 99832 30436 99888 30492
rect 99888 30436 99892 30492
rect 99828 30432 99892 30436
rect 99908 30492 99972 30496
rect 99908 30436 99912 30492
rect 99912 30436 99968 30492
rect 99968 30436 99972 30492
rect 99908 30432 99972 30436
rect 1308 29948 1372 29952
rect 1308 29892 1312 29948
rect 1312 29892 1368 29948
rect 1368 29892 1372 29948
rect 1308 29888 1372 29892
rect 1388 29948 1452 29952
rect 1388 29892 1392 29948
rect 1392 29892 1448 29948
rect 1448 29892 1452 29948
rect 1388 29888 1452 29892
rect 98932 29948 98996 29952
rect 98932 29892 98936 29948
rect 98936 29892 98992 29948
rect 98992 29892 98996 29948
rect 98932 29888 98996 29892
rect 99012 29948 99076 29952
rect 99012 29892 99016 29948
rect 99016 29892 99072 29948
rect 99072 29892 99076 29948
rect 99012 29888 99076 29892
rect 99092 29948 99156 29952
rect 99092 29892 99096 29948
rect 99096 29892 99152 29948
rect 99152 29892 99156 29948
rect 99092 29888 99156 29892
rect 99172 29948 99236 29952
rect 99172 29892 99176 29948
rect 99176 29892 99232 29948
rect 99232 29892 99236 29948
rect 99172 29888 99236 29892
rect 1676 29404 1740 29408
rect 1676 29348 1680 29404
rect 1680 29348 1736 29404
rect 1736 29348 1740 29404
rect 1676 29344 1740 29348
rect 1756 29404 1820 29408
rect 1756 29348 1760 29404
rect 1760 29348 1816 29404
rect 1816 29348 1820 29404
rect 1756 29344 1820 29348
rect 99668 29404 99732 29408
rect 99668 29348 99672 29404
rect 99672 29348 99728 29404
rect 99728 29348 99732 29404
rect 99668 29344 99732 29348
rect 99748 29404 99812 29408
rect 99748 29348 99752 29404
rect 99752 29348 99808 29404
rect 99808 29348 99812 29404
rect 99748 29344 99812 29348
rect 99828 29404 99892 29408
rect 99828 29348 99832 29404
rect 99832 29348 99888 29404
rect 99888 29348 99892 29404
rect 99828 29344 99892 29348
rect 99908 29404 99972 29408
rect 99908 29348 99912 29404
rect 99912 29348 99968 29404
rect 99968 29348 99972 29404
rect 99908 29344 99972 29348
rect 1308 28860 1372 28864
rect 1308 28804 1312 28860
rect 1312 28804 1368 28860
rect 1368 28804 1372 28860
rect 1308 28800 1372 28804
rect 1388 28860 1452 28864
rect 1388 28804 1392 28860
rect 1392 28804 1448 28860
rect 1448 28804 1452 28860
rect 1388 28800 1452 28804
rect 98932 28860 98996 28864
rect 98932 28804 98936 28860
rect 98936 28804 98992 28860
rect 98992 28804 98996 28860
rect 98932 28800 98996 28804
rect 99012 28860 99076 28864
rect 99012 28804 99016 28860
rect 99016 28804 99072 28860
rect 99072 28804 99076 28860
rect 99012 28800 99076 28804
rect 99092 28860 99156 28864
rect 99092 28804 99096 28860
rect 99096 28804 99152 28860
rect 99152 28804 99156 28860
rect 99092 28800 99156 28804
rect 99172 28860 99236 28864
rect 99172 28804 99176 28860
rect 99176 28804 99232 28860
rect 99232 28804 99236 28860
rect 99172 28800 99236 28804
rect 1676 28316 1740 28320
rect 1676 28260 1680 28316
rect 1680 28260 1736 28316
rect 1736 28260 1740 28316
rect 1676 28256 1740 28260
rect 1756 28316 1820 28320
rect 1756 28260 1760 28316
rect 1760 28260 1816 28316
rect 1816 28260 1820 28316
rect 1756 28256 1820 28260
rect 99668 28316 99732 28320
rect 99668 28260 99672 28316
rect 99672 28260 99728 28316
rect 99728 28260 99732 28316
rect 99668 28256 99732 28260
rect 99748 28316 99812 28320
rect 99748 28260 99752 28316
rect 99752 28260 99808 28316
rect 99808 28260 99812 28316
rect 99748 28256 99812 28260
rect 99828 28316 99892 28320
rect 99828 28260 99832 28316
rect 99832 28260 99888 28316
rect 99888 28260 99892 28316
rect 99828 28256 99892 28260
rect 99908 28316 99972 28320
rect 99908 28260 99912 28316
rect 99912 28260 99968 28316
rect 99968 28260 99972 28316
rect 99908 28256 99972 28260
rect 1308 27772 1372 27776
rect 1308 27716 1312 27772
rect 1312 27716 1368 27772
rect 1368 27716 1372 27772
rect 1308 27712 1372 27716
rect 1388 27772 1452 27776
rect 1388 27716 1392 27772
rect 1392 27716 1448 27772
rect 1448 27716 1452 27772
rect 1388 27712 1452 27716
rect 98932 27772 98996 27776
rect 98932 27716 98936 27772
rect 98936 27716 98992 27772
rect 98992 27716 98996 27772
rect 98932 27712 98996 27716
rect 99012 27772 99076 27776
rect 99012 27716 99016 27772
rect 99016 27716 99072 27772
rect 99072 27716 99076 27772
rect 99012 27712 99076 27716
rect 99092 27772 99156 27776
rect 99092 27716 99096 27772
rect 99096 27716 99152 27772
rect 99152 27716 99156 27772
rect 99092 27712 99156 27716
rect 99172 27772 99236 27776
rect 99172 27716 99176 27772
rect 99176 27716 99232 27772
rect 99232 27716 99236 27772
rect 99172 27712 99236 27716
rect 1676 27228 1740 27232
rect 1676 27172 1680 27228
rect 1680 27172 1736 27228
rect 1736 27172 1740 27228
rect 1676 27168 1740 27172
rect 1756 27228 1820 27232
rect 1756 27172 1760 27228
rect 1760 27172 1816 27228
rect 1816 27172 1820 27228
rect 1756 27168 1820 27172
rect 99668 27228 99732 27232
rect 99668 27172 99672 27228
rect 99672 27172 99728 27228
rect 99728 27172 99732 27228
rect 99668 27168 99732 27172
rect 99748 27228 99812 27232
rect 99748 27172 99752 27228
rect 99752 27172 99808 27228
rect 99808 27172 99812 27228
rect 99748 27168 99812 27172
rect 99828 27228 99892 27232
rect 99828 27172 99832 27228
rect 99832 27172 99888 27228
rect 99888 27172 99892 27228
rect 99828 27168 99892 27172
rect 99908 27228 99972 27232
rect 99908 27172 99912 27228
rect 99912 27172 99968 27228
rect 99968 27172 99972 27228
rect 99908 27168 99972 27172
rect 1308 26684 1372 26688
rect 1308 26628 1312 26684
rect 1312 26628 1368 26684
rect 1368 26628 1372 26684
rect 1308 26624 1372 26628
rect 1388 26684 1452 26688
rect 1388 26628 1392 26684
rect 1392 26628 1448 26684
rect 1448 26628 1452 26684
rect 1388 26624 1452 26628
rect 98932 26684 98996 26688
rect 98932 26628 98936 26684
rect 98936 26628 98992 26684
rect 98992 26628 98996 26684
rect 98932 26624 98996 26628
rect 99012 26684 99076 26688
rect 99012 26628 99016 26684
rect 99016 26628 99072 26684
rect 99072 26628 99076 26684
rect 99012 26624 99076 26628
rect 99092 26684 99156 26688
rect 99092 26628 99096 26684
rect 99096 26628 99152 26684
rect 99152 26628 99156 26684
rect 99092 26624 99156 26628
rect 99172 26684 99236 26688
rect 99172 26628 99176 26684
rect 99176 26628 99232 26684
rect 99232 26628 99236 26684
rect 99172 26624 99236 26628
rect 1676 26140 1740 26144
rect 1676 26084 1680 26140
rect 1680 26084 1736 26140
rect 1736 26084 1740 26140
rect 1676 26080 1740 26084
rect 1756 26140 1820 26144
rect 1756 26084 1760 26140
rect 1760 26084 1816 26140
rect 1816 26084 1820 26140
rect 1756 26080 1820 26084
rect 99668 26140 99732 26144
rect 99668 26084 99672 26140
rect 99672 26084 99728 26140
rect 99728 26084 99732 26140
rect 99668 26080 99732 26084
rect 99748 26140 99812 26144
rect 99748 26084 99752 26140
rect 99752 26084 99808 26140
rect 99808 26084 99812 26140
rect 99748 26080 99812 26084
rect 99828 26140 99892 26144
rect 99828 26084 99832 26140
rect 99832 26084 99888 26140
rect 99888 26084 99892 26140
rect 99828 26080 99892 26084
rect 99908 26140 99972 26144
rect 99908 26084 99912 26140
rect 99912 26084 99968 26140
rect 99968 26084 99972 26140
rect 99908 26080 99972 26084
rect 1308 25596 1372 25600
rect 1308 25540 1312 25596
rect 1312 25540 1368 25596
rect 1368 25540 1372 25596
rect 1308 25536 1372 25540
rect 1388 25596 1452 25600
rect 1388 25540 1392 25596
rect 1392 25540 1448 25596
rect 1448 25540 1452 25596
rect 1388 25536 1452 25540
rect 98932 25596 98996 25600
rect 98932 25540 98936 25596
rect 98936 25540 98992 25596
rect 98992 25540 98996 25596
rect 98932 25536 98996 25540
rect 99012 25596 99076 25600
rect 99012 25540 99016 25596
rect 99016 25540 99072 25596
rect 99072 25540 99076 25596
rect 99012 25536 99076 25540
rect 99092 25596 99156 25600
rect 99092 25540 99096 25596
rect 99096 25540 99152 25596
rect 99152 25540 99156 25596
rect 99092 25536 99156 25540
rect 99172 25596 99236 25600
rect 99172 25540 99176 25596
rect 99176 25540 99232 25596
rect 99232 25540 99236 25596
rect 99172 25536 99236 25540
rect 1676 25052 1740 25056
rect 1676 24996 1680 25052
rect 1680 24996 1736 25052
rect 1736 24996 1740 25052
rect 1676 24992 1740 24996
rect 1756 25052 1820 25056
rect 1756 24996 1760 25052
rect 1760 24996 1816 25052
rect 1816 24996 1820 25052
rect 1756 24992 1820 24996
rect 99668 25052 99732 25056
rect 99668 24996 99672 25052
rect 99672 24996 99728 25052
rect 99728 24996 99732 25052
rect 99668 24992 99732 24996
rect 99748 25052 99812 25056
rect 99748 24996 99752 25052
rect 99752 24996 99808 25052
rect 99808 24996 99812 25052
rect 99748 24992 99812 24996
rect 99828 25052 99892 25056
rect 99828 24996 99832 25052
rect 99832 24996 99888 25052
rect 99888 24996 99892 25052
rect 99828 24992 99892 24996
rect 99908 25052 99972 25056
rect 99908 24996 99912 25052
rect 99912 24996 99968 25052
rect 99968 24996 99972 25052
rect 99908 24992 99972 24996
rect 1308 24508 1372 24512
rect 1308 24452 1312 24508
rect 1312 24452 1368 24508
rect 1368 24452 1372 24508
rect 1308 24448 1372 24452
rect 1388 24508 1452 24512
rect 1388 24452 1392 24508
rect 1392 24452 1448 24508
rect 1448 24452 1452 24508
rect 1388 24448 1452 24452
rect 98932 24508 98996 24512
rect 98932 24452 98936 24508
rect 98936 24452 98992 24508
rect 98992 24452 98996 24508
rect 98932 24448 98996 24452
rect 99012 24508 99076 24512
rect 99012 24452 99016 24508
rect 99016 24452 99072 24508
rect 99072 24452 99076 24508
rect 99012 24448 99076 24452
rect 99092 24508 99156 24512
rect 99092 24452 99096 24508
rect 99096 24452 99152 24508
rect 99152 24452 99156 24508
rect 99092 24448 99156 24452
rect 99172 24508 99236 24512
rect 99172 24452 99176 24508
rect 99176 24452 99232 24508
rect 99232 24452 99236 24508
rect 99172 24448 99236 24452
rect 1676 23964 1740 23968
rect 1676 23908 1680 23964
rect 1680 23908 1736 23964
rect 1736 23908 1740 23964
rect 1676 23904 1740 23908
rect 1756 23964 1820 23968
rect 1756 23908 1760 23964
rect 1760 23908 1816 23964
rect 1816 23908 1820 23964
rect 1756 23904 1820 23908
rect 99668 23964 99732 23968
rect 99668 23908 99672 23964
rect 99672 23908 99728 23964
rect 99728 23908 99732 23964
rect 99668 23904 99732 23908
rect 99748 23964 99812 23968
rect 99748 23908 99752 23964
rect 99752 23908 99808 23964
rect 99808 23908 99812 23964
rect 99748 23904 99812 23908
rect 99828 23964 99892 23968
rect 99828 23908 99832 23964
rect 99832 23908 99888 23964
rect 99888 23908 99892 23964
rect 99828 23904 99892 23908
rect 99908 23964 99972 23968
rect 99908 23908 99912 23964
rect 99912 23908 99968 23964
rect 99968 23908 99972 23964
rect 99908 23904 99972 23908
rect 1308 23420 1372 23424
rect 1308 23364 1312 23420
rect 1312 23364 1368 23420
rect 1368 23364 1372 23420
rect 1308 23360 1372 23364
rect 1388 23420 1452 23424
rect 1388 23364 1392 23420
rect 1392 23364 1448 23420
rect 1448 23364 1452 23420
rect 1388 23360 1452 23364
rect 98932 23420 98996 23424
rect 98932 23364 98936 23420
rect 98936 23364 98992 23420
rect 98992 23364 98996 23420
rect 98932 23360 98996 23364
rect 99012 23420 99076 23424
rect 99012 23364 99016 23420
rect 99016 23364 99072 23420
rect 99072 23364 99076 23420
rect 99012 23360 99076 23364
rect 99092 23420 99156 23424
rect 99092 23364 99096 23420
rect 99096 23364 99152 23420
rect 99152 23364 99156 23420
rect 99092 23360 99156 23364
rect 99172 23420 99236 23424
rect 99172 23364 99176 23420
rect 99176 23364 99232 23420
rect 99232 23364 99236 23420
rect 99172 23360 99236 23364
rect 1676 22876 1740 22880
rect 1676 22820 1680 22876
rect 1680 22820 1736 22876
rect 1736 22820 1740 22876
rect 1676 22816 1740 22820
rect 1756 22876 1820 22880
rect 1756 22820 1760 22876
rect 1760 22820 1816 22876
rect 1816 22820 1820 22876
rect 1756 22816 1820 22820
rect 99668 22876 99732 22880
rect 99668 22820 99672 22876
rect 99672 22820 99728 22876
rect 99728 22820 99732 22876
rect 99668 22816 99732 22820
rect 99748 22876 99812 22880
rect 99748 22820 99752 22876
rect 99752 22820 99808 22876
rect 99808 22820 99812 22876
rect 99748 22816 99812 22820
rect 99828 22876 99892 22880
rect 99828 22820 99832 22876
rect 99832 22820 99888 22876
rect 99888 22820 99892 22876
rect 99828 22816 99892 22820
rect 99908 22876 99972 22880
rect 99908 22820 99912 22876
rect 99912 22820 99968 22876
rect 99968 22820 99972 22876
rect 99908 22816 99972 22820
rect 1308 22332 1372 22336
rect 1308 22276 1312 22332
rect 1312 22276 1368 22332
rect 1368 22276 1372 22332
rect 1308 22272 1372 22276
rect 1388 22332 1452 22336
rect 1388 22276 1392 22332
rect 1392 22276 1448 22332
rect 1448 22276 1452 22332
rect 1388 22272 1452 22276
rect 98932 22332 98996 22336
rect 98932 22276 98936 22332
rect 98936 22276 98992 22332
rect 98992 22276 98996 22332
rect 98932 22272 98996 22276
rect 99012 22332 99076 22336
rect 99012 22276 99016 22332
rect 99016 22276 99072 22332
rect 99072 22276 99076 22332
rect 99012 22272 99076 22276
rect 99092 22332 99156 22336
rect 99092 22276 99096 22332
rect 99096 22276 99152 22332
rect 99152 22276 99156 22332
rect 99092 22272 99156 22276
rect 99172 22332 99236 22336
rect 99172 22276 99176 22332
rect 99176 22276 99232 22332
rect 99232 22276 99236 22332
rect 99172 22272 99236 22276
rect 1676 21788 1740 21792
rect 1676 21732 1680 21788
rect 1680 21732 1736 21788
rect 1736 21732 1740 21788
rect 1676 21728 1740 21732
rect 1756 21788 1820 21792
rect 1756 21732 1760 21788
rect 1760 21732 1816 21788
rect 1816 21732 1820 21788
rect 1756 21728 1820 21732
rect 99668 21788 99732 21792
rect 99668 21732 99672 21788
rect 99672 21732 99728 21788
rect 99728 21732 99732 21788
rect 99668 21728 99732 21732
rect 99748 21788 99812 21792
rect 99748 21732 99752 21788
rect 99752 21732 99808 21788
rect 99808 21732 99812 21788
rect 99748 21728 99812 21732
rect 99828 21788 99892 21792
rect 99828 21732 99832 21788
rect 99832 21732 99888 21788
rect 99888 21732 99892 21788
rect 99828 21728 99892 21732
rect 99908 21788 99972 21792
rect 99908 21732 99912 21788
rect 99912 21732 99968 21788
rect 99968 21732 99972 21788
rect 99908 21728 99972 21732
rect 1308 21244 1372 21248
rect 1308 21188 1312 21244
rect 1312 21188 1368 21244
rect 1368 21188 1372 21244
rect 1308 21184 1372 21188
rect 1388 21244 1452 21248
rect 1388 21188 1392 21244
rect 1392 21188 1448 21244
rect 1448 21188 1452 21244
rect 1388 21184 1452 21188
rect 98932 21244 98996 21248
rect 98932 21188 98936 21244
rect 98936 21188 98992 21244
rect 98992 21188 98996 21244
rect 98932 21184 98996 21188
rect 99012 21244 99076 21248
rect 99012 21188 99016 21244
rect 99016 21188 99072 21244
rect 99072 21188 99076 21244
rect 99012 21184 99076 21188
rect 99092 21244 99156 21248
rect 99092 21188 99096 21244
rect 99096 21188 99152 21244
rect 99152 21188 99156 21244
rect 99092 21184 99156 21188
rect 99172 21244 99236 21248
rect 99172 21188 99176 21244
rect 99176 21188 99232 21244
rect 99232 21188 99236 21244
rect 99172 21184 99236 21188
rect 1676 20700 1740 20704
rect 1676 20644 1680 20700
rect 1680 20644 1736 20700
rect 1736 20644 1740 20700
rect 1676 20640 1740 20644
rect 1756 20700 1820 20704
rect 1756 20644 1760 20700
rect 1760 20644 1816 20700
rect 1816 20644 1820 20700
rect 1756 20640 1820 20644
rect 99668 20700 99732 20704
rect 99668 20644 99672 20700
rect 99672 20644 99728 20700
rect 99728 20644 99732 20700
rect 99668 20640 99732 20644
rect 99748 20700 99812 20704
rect 99748 20644 99752 20700
rect 99752 20644 99808 20700
rect 99808 20644 99812 20700
rect 99748 20640 99812 20644
rect 99828 20700 99892 20704
rect 99828 20644 99832 20700
rect 99832 20644 99888 20700
rect 99888 20644 99892 20700
rect 99828 20640 99892 20644
rect 99908 20700 99972 20704
rect 99908 20644 99912 20700
rect 99912 20644 99968 20700
rect 99968 20644 99972 20700
rect 99908 20640 99972 20644
rect 1308 20156 1372 20160
rect 1308 20100 1312 20156
rect 1312 20100 1368 20156
rect 1368 20100 1372 20156
rect 1308 20096 1372 20100
rect 1388 20156 1452 20160
rect 1388 20100 1392 20156
rect 1392 20100 1448 20156
rect 1448 20100 1452 20156
rect 1388 20096 1452 20100
rect 98932 20156 98996 20160
rect 98932 20100 98936 20156
rect 98936 20100 98992 20156
rect 98992 20100 98996 20156
rect 98932 20096 98996 20100
rect 99012 20156 99076 20160
rect 99012 20100 99016 20156
rect 99016 20100 99072 20156
rect 99072 20100 99076 20156
rect 99012 20096 99076 20100
rect 99092 20156 99156 20160
rect 99092 20100 99096 20156
rect 99096 20100 99152 20156
rect 99152 20100 99156 20156
rect 99092 20096 99156 20100
rect 99172 20156 99236 20160
rect 99172 20100 99176 20156
rect 99176 20100 99232 20156
rect 99232 20100 99236 20156
rect 99172 20096 99236 20100
rect 1676 19612 1740 19616
rect 1676 19556 1680 19612
rect 1680 19556 1736 19612
rect 1736 19556 1740 19612
rect 1676 19552 1740 19556
rect 1756 19612 1820 19616
rect 1756 19556 1760 19612
rect 1760 19556 1816 19612
rect 1816 19556 1820 19612
rect 1756 19552 1820 19556
rect 99668 19612 99732 19616
rect 99668 19556 99672 19612
rect 99672 19556 99728 19612
rect 99728 19556 99732 19612
rect 99668 19552 99732 19556
rect 99748 19612 99812 19616
rect 99748 19556 99752 19612
rect 99752 19556 99808 19612
rect 99808 19556 99812 19612
rect 99748 19552 99812 19556
rect 99828 19612 99892 19616
rect 99828 19556 99832 19612
rect 99832 19556 99888 19612
rect 99888 19556 99892 19612
rect 99828 19552 99892 19556
rect 99908 19612 99972 19616
rect 99908 19556 99912 19612
rect 99912 19556 99968 19612
rect 99968 19556 99972 19612
rect 99908 19552 99972 19556
rect 1308 19068 1372 19072
rect 1308 19012 1312 19068
rect 1312 19012 1368 19068
rect 1368 19012 1372 19068
rect 1308 19008 1372 19012
rect 1388 19068 1452 19072
rect 1388 19012 1392 19068
rect 1392 19012 1448 19068
rect 1448 19012 1452 19068
rect 1388 19008 1452 19012
rect 98932 19068 98996 19072
rect 98932 19012 98936 19068
rect 98936 19012 98992 19068
rect 98992 19012 98996 19068
rect 98932 19008 98996 19012
rect 99012 19068 99076 19072
rect 99012 19012 99016 19068
rect 99016 19012 99072 19068
rect 99072 19012 99076 19068
rect 99012 19008 99076 19012
rect 99092 19068 99156 19072
rect 99092 19012 99096 19068
rect 99096 19012 99152 19068
rect 99152 19012 99156 19068
rect 99092 19008 99156 19012
rect 99172 19068 99236 19072
rect 99172 19012 99176 19068
rect 99176 19012 99232 19068
rect 99232 19012 99236 19068
rect 99172 19008 99236 19012
rect 1676 18524 1740 18528
rect 1676 18468 1680 18524
rect 1680 18468 1736 18524
rect 1736 18468 1740 18524
rect 1676 18464 1740 18468
rect 1756 18524 1820 18528
rect 1756 18468 1760 18524
rect 1760 18468 1816 18524
rect 1816 18468 1820 18524
rect 1756 18464 1820 18468
rect 99668 18524 99732 18528
rect 99668 18468 99672 18524
rect 99672 18468 99728 18524
rect 99728 18468 99732 18524
rect 99668 18464 99732 18468
rect 99748 18524 99812 18528
rect 99748 18468 99752 18524
rect 99752 18468 99808 18524
rect 99808 18468 99812 18524
rect 99748 18464 99812 18468
rect 99828 18524 99892 18528
rect 99828 18468 99832 18524
rect 99832 18468 99888 18524
rect 99888 18468 99892 18524
rect 99828 18464 99892 18468
rect 99908 18524 99972 18528
rect 99908 18468 99912 18524
rect 99912 18468 99968 18524
rect 99968 18468 99972 18524
rect 99908 18464 99972 18468
rect 1308 17980 1372 17984
rect 1308 17924 1312 17980
rect 1312 17924 1368 17980
rect 1368 17924 1372 17980
rect 1308 17920 1372 17924
rect 1388 17980 1452 17984
rect 1388 17924 1392 17980
rect 1392 17924 1448 17980
rect 1448 17924 1452 17980
rect 1388 17920 1452 17924
rect 98932 17980 98996 17984
rect 98932 17924 98936 17980
rect 98936 17924 98992 17980
rect 98992 17924 98996 17980
rect 98932 17920 98996 17924
rect 99012 17980 99076 17984
rect 99012 17924 99016 17980
rect 99016 17924 99072 17980
rect 99072 17924 99076 17980
rect 99012 17920 99076 17924
rect 99092 17980 99156 17984
rect 99092 17924 99096 17980
rect 99096 17924 99152 17980
rect 99152 17924 99156 17980
rect 99092 17920 99156 17924
rect 99172 17980 99236 17984
rect 99172 17924 99176 17980
rect 99176 17924 99232 17980
rect 99232 17924 99236 17980
rect 99172 17920 99236 17924
rect 1676 17436 1740 17440
rect 1676 17380 1680 17436
rect 1680 17380 1736 17436
rect 1736 17380 1740 17436
rect 1676 17376 1740 17380
rect 1756 17436 1820 17440
rect 1756 17380 1760 17436
rect 1760 17380 1816 17436
rect 1816 17380 1820 17436
rect 1756 17376 1820 17380
rect 99668 17436 99732 17440
rect 99668 17380 99672 17436
rect 99672 17380 99728 17436
rect 99728 17380 99732 17436
rect 99668 17376 99732 17380
rect 99748 17436 99812 17440
rect 99748 17380 99752 17436
rect 99752 17380 99808 17436
rect 99808 17380 99812 17436
rect 99748 17376 99812 17380
rect 99828 17436 99892 17440
rect 99828 17380 99832 17436
rect 99832 17380 99888 17436
rect 99888 17380 99892 17436
rect 99828 17376 99892 17380
rect 99908 17436 99972 17440
rect 99908 17380 99912 17436
rect 99912 17380 99968 17436
rect 99968 17380 99972 17436
rect 99908 17376 99972 17380
rect 1308 16892 1372 16896
rect 1308 16836 1312 16892
rect 1312 16836 1368 16892
rect 1368 16836 1372 16892
rect 1308 16832 1372 16836
rect 1388 16892 1452 16896
rect 1388 16836 1392 16892
rect 1392 16836 1448 16892
rect 1448 16836 1452 16892
rect 1388 16832 1452 16836
rect 98932 16892 98996 16896
rect 98932 16836 98936 16892
rect 98936 16836 98992 16892
rect 98992 16836 98996 16892
rect 98932 16832 98996 16836
rect 99012 16892 99076 16896
rect 99012 16836 99016 16892
rect 99016 16836 99072 16892
rect 99072 16836 99076 16892
rect 99012 16832 99076 16836
rect 99092 16892 99156 16896
rect 99092 16836 99096 16892
rect 99096 16836 99152 16892
rect 99152 16836 99156 16892
rect 99092 16832 99156 16836
rect 99172 16892 99236 16896
rect 99172 16836 99176 16892
rect 99176 16836 99232 16892
rect 99232 16836 99236 16892
rect 99172 16832 99236 16836
rect 1676 16348 1740 16352
rect 1676 16292 1680 16348
rect 1680 16292 1736 16348
rect 1736 16292 1740 16348
rect 1676 16288 1740 16292
rect 1756 16348 1820 16352
rect 1756 16292 1760 16348
rect 1760 16292 1816 16348
rect 1816 16292 1820 16348
rect 1756 16288 1820 16292
rect 99668 16348 99732 16352
rect 99668 16292 99672 16348
rect 99672 16292 99728 16348
rect 99728 16292 99732 16348
rect 99668 16288 99732 16292
rect 99748 16348 99812 16352
rect 99748 16292 99752 16348
rect 99752 16292 99808 16348
rect 99808 16292 99812 16348
rect 99748 16288 99812 16292
rect 99828 16348 99892 16352
rect 99828 16292 99832 16348
rect 99832 16292 99888 16348
rect 99888 16292 99892 16348
rect 99828 16288 99892 16292
rect 99908 16348 99972 16352
rect 99908 16292 99912 16348
rect 99912 16292 99968 16348
rect 99968 16292 99972 16348
rect 99908 16288 99972 16292
rect 1308 15804 1372 15808
rect 1308 15748 1312 15804
rect 1312 15748 1368 15804
rect 1368 15748 1372 15804
rect 1308 15744 1372 15748
rect 1388 15804 1452 15808
rect 1388 15748 1392 15804
rect 1392 15748 1448 15804
rect 1448 15748 1452 15804
rect 1388 15744 1452 15748
rect 98932 15804 98996 15808
rect 98932 15748 98936 15804
rect 98936 15748 98992 15804
rect 98992 15748 98996 15804
rect 98932 15744 98996 15748
rect 99012 15804 99076 15808
rect 99012 15748 99016 15804
rect 99016 15748 99072 15804
rect 99072 15748 99076 15804
rect 99012 15744 99076 15748
rect 99092 15804 99156 15808
rect 99092 15748 99096 15804
rect 99096 15748 99152 15804
rect 99152 15748 99156 15804
rect 99092 15744 99156 15748
rect 99172 15804 99236 15808
rect 99172 15748 99176 15804
rect 99176 15748 99232 15804
rect 99232 15748 99236 15804
rect 99172 15744 99236 15748
rect 1676 15260 1740 15264
rect 1676 15204 1680 15260
rect 1680 15204 1736 15260
rect 1736 15204 1740 15260
rect 1676 15200 1740 15204
rect 1756 15260 1820 15264
rect 1756 15204 1760 15260
rect 1760 15204 1816 15260
rect 1816 15204 1820 15260
rect 1756 15200 1820 15204
rect 99668 15260 99732 15264
rect 99668 15204 99672 15260
rect 99672 15204 99728 15260
rect 99728 15204 99732 15260
rect 99668 15200 99732 15204
rect 99748 15260 99812 15264
rect 99748 15204 99752 15260
rect 99752 15204 99808 15260
rect 99808 15204 99812 15260
rect 99748 15200 99812 15204
rect 99828 15260 99892 15264
rect 99828 15204 99832 15260
rect 99832 15204 99888 15260
rect 99888 15204 99892 15260
rect 99828 15200 99892 15204
rect 99908 15260 99972 15264
rect 99908 15204 99912 15260
rect 99912 15204 99968 15260
rect 99968 15204 99972 15260
rect 99908 15200 99972 15204
rect 1308 14716 1372 14720
rect 1308 14660 1312 14716
rect 1312 14660 1368 14716
rect 1368 14660 1372 14716
rect 1308 14656 1372 14660
rect 1388 14716 1452 14720
rect 1388 14660 1392 14716
rect 1392 14660 1448 14716
rect 1448 14660 1452 14716
rect 1388 14656 1452 14660
rect 98932 14716 98996 14720
rect 98932 14660 98936 14716
rect 98936 14660 98992 14716
rect 98992 14660 98996 14716
rect 98932 14656 98996 14660
rect 99012 14716 99076 14720
rect 99012 14660 99016 14716
rect 99016 14660 99072 14716
rect 99072 14660 99076 14716
rect 99012 14656 99076 14660
rect 99092 14716 99156 14720
rect 99092 14660 99096 14716
rect 99096 14660 99152 14716
rect 99152 14660 99156 14716
rect 99092 14656 99156 14660
rect 99172 14716 99236 14720
rect 99172 14660 99176 14716
rect 99176 14660 99232 14716
rect 99232 14660 99236 14716
rect 99172 14656 99236 14660
rect 1676 14172 1740 14176
rect 1676 14116 1680 14172
rect 1680 14116 1736 14172
rect 1736 14116 1740 14172
rect 1676 14112 1740 14116
rect 1756 14172 1820 14176
rect 1756 14116 1760 14172
rect 1760 14116 1816 14172
rect 1816 14116 1820 14172
rect 1756 14112 1820 14116
rect 99668 14172 99732 14176
rect 99668 14116 99672 14172
rect 99672 14116 99728 14172
rect 99728 14116 99732 14172
rect 99668 14112 99732 14116
rect 99748 14172 99812 14176
rect 99748 14116 99752 14172
rect 99752 14116 99808 14172
rect 99808 14116 99812 14172
rect 99748 14112 99812 14116
rect 99828 14172 99892 14176
rect 99828 14116 99832 14172
rect 99832 14116 99888 14172
rect 99888 14116 99892 14172
rect 99828 14112 99892 14116
rect 99908 14172 99972 14176
rect 99908 14116 99912 14172
rect 99912 14116 99968 14172
rect 99968 14116 99972 14172
rect 99908 14112 99972 14116
rect 1308 13628 1372 13632
rect 1308 13572 1312 13628
rect 1312 13572 1368 13628
rect 1368 13572 1372 13628
rect 1308 13568 1372 13572
rect 1388 13628 1452 13632
rect 1388 13572 1392 13628
rect 1392 13572 1448 13628
rect 1448 13572 1452 13628
rect 1388 13568 1452 13572
rect 98932 13628 98996 13632
rect 98932 13572 98936 13628
rect 98936 13572 98992 13628
rect 98992 13572 98996 13628
rect 98932 13568 98996 13572
rect 99012 13628 99076 13632
rect 99012 13572 99016 13628
rect 99016 13572 99072 13628
rect 99072 13572 99076 13628
rect 99012 13568 99076 13572
rect 99092 13628 99156 13632
rect 99092 13572 99096 13628
rect 99096 13572 99152 13628
rect 99152 13572 99156 13628
rect 99092 13568 99156 13572
rect 99172 13628 99236 13632
rect 99172 13572 99176 13628
rect 99176 13572 99232 13628
rect 99232 13572 99236 13628
rect 99172 13568 99236 13572
rect 1676 13084 1740 13088
rect 1676 13028 1680 13084
rect 1680 13028 1736 13084
rect 1736 13028 1740 13084
rect 1676 13024 1740 13028
rect 1756 13084 1820 13088
rect 1756 13028 1760 13084
rect 1760 13028 1816 13084
rect 1816 13028 1820 13084
rect 1756 13024 1820 13028
rect 99668 13084 99732 13088
rect 99668 13028 99672 13084
rect 99672 13028 99728 13084
rect 99728 13028 99732 13084
rect 99668 13024 99732 13028
rect 99748 13084 99812 13088
rect 99748 13028 99752 13084
rect 99752 13028 99808 13084
rect 99808 13028 99812 13084
rect 99748 13024 99812 13028
rect 99828 13084 99892 13088
rect 99828 13028 99832 13084
rect 99832 13028 99888 13084
rect 99888 13028 99892 13084
rect 99828 13024 99892 13028
rect 99908 13084 99972 13088
rect 99908 13028 99912 13084
rect 99912 13028 99968 13084
rect 99968 13028 99972 13084
rect 99908 13024 99972 13028
rect 1308 12540 1372 12544
rect 1308 12484 1312 12540
rect 1312 12484 1368 12540
rect 1368 12484 1372 12540
rect 1308 12480 1372 12484
rect 1388 12540 1452 12544
rect 1388 12484 1392 12540
rect 1392 12484 1448 12540
rect 1448 12484 1452 12540
rect 1388 12480 1452 12484
rect 98932 12540 98996 12544
rect 98932 12484 98936 12540
rect 98936 12484 98992 12540
rect 98992 12484 98996 12540
rect 98932 12480 98996 12484
rect 99012 12540 99076 12544
rect 99012 12484 99016 12540
rect 99016 12484 99072 12540
rect 99072 12484 99076 12540
rect 99012 12480 99076 12484
rect 99092 12540 99156 12544
rect 99092 12484 99096 12540
rect 99096 12484 99152 12540
rect 99152 12484 99156 12540
rect 99092 12480 99156 12484
rect 99172 12540 99236 12544
rect 99172 12484 99176 12540
rect 99176 12484 99232 12540
rect 99232 12484 99236 12540
rect 99172 12480 99236 12484
rect 1676 11996 1740 12000
rect 1676 11940 1680 11996
rect 1680 11940 1736 11996
rect 1736 11940 1740 11996
rect 1676 11936 1740 11940
rect 1756 11996 1820 12000
rect 1756 11940 1760 11996
rect 1760 11940 1816 11996
rect 1816 11940 1820 11996
rect 1756 11936 1820 11940
rect 99668 11996 99732 12000
rect 99668 11940 99672 11996
rect 99672 11940 99728 11996
rect 99728 11940 99732 11996
rect 99668 11936 99732 11940
rect 99748 11996 99812 12000
rect 99748 11940 99752 11996
rect 99752 11940 99808 11996
rect 99808 11940 99812 11996
rect 99748 11936 99812 11940
rect 99828 11996 99892 12000
rect 99828 11940 99832 11996
rect 99832 11940 99888 11996
rect 99888 11940 99892 11996
rect 99828 11936 99892 11940
rect 99908 11996 99972 12000
rect 99908 11940 99912 11996
rect 99912 11940 99968 11996
rect 99968 11940 99972 11996
rect 99908 11936 99972 11940
rect 1308 11452 1372 11456
rect 1308 11396 1312 11452
rect 1312 11396 1368 11452
rect 1368 11396 1372 11452
rect 1308 11392 1372 11396
rect 1388 11452 1452 11456
rect 1388 11396 1392 11452
rect 1392 11396 1448 11452
rect 1448 11396 1452 11452
rect 1388 11392 1452 11396
rect 98932 11452 98996 11456
rect 98932 11396 98936 11452
rect 98936 11396 98992 11452
rect 98992 11396 98996 11452
rect 98932 11392 98996 11396
rect 99012 11452 99076 11456
rect 99012 11396 99016 11452
rect 99016 11396 99072 11452
rect 99072 11396 99076 11452
rect 99012 11392 99076 11396
rect 99092 11452 99156 11456
rect 99092 11396 99096 11452
rect 99096 11396 99152 11452
rect 99152 11396 99156 11452
rect 99092 11392 99156 11396
rect 99172 11452 99236 11456
rect 99172 11396 99176 11452
rect 99176 11396 99232 11452
rect 99232 11396 99236 11452
rect 99172 11392 99236 11396
rect 1676 10908 1740 10912
rect 1676 10852 1680 10908
rect 1680 10852 1736 10908
rect 1736 10852 1740 10908
rect 1676 10848 1740 10852
rect 1756 10908 1820 10912
rect 1756 10852 1760 10908
rect 1760 10852 1816 10908
rect 1816 10852 1820 10908
rect 1756 10848 1820 10852
rect 99668 10908 99732 10912
rect 99668 10852 99672 10908
rect 99672 10852 99728 10908
rect 99728 10852 99732 10908
rect 99668 10848 99732 10852
rect 99748 10908 99812 10912
rect 99748 10852 99752 10908
rect 99752 10852 99808 10908
rect 99808 10852 99812 10908
rect 99748 10848 99812 10852
rect 99828 10908 99892 10912
rect 99828 10852 99832 10908
rect 99832 10852 99888 10908
rect 99888 10852 99892 10908
rect 99828 10848 99892 10852
rect 99908 10908 99972 10912
rect 99908 10852 99912 10908
rect 99912 10852 99968 10908
rect 99968 10852 99972 10908
rect 99908 10848 99972 10852
rect 1308 10364 1372 10368
rect 1308 10308 1312 10364
rect 1312 10308 1368 10364
rect 1368 10308 1372 10364
rect 1308 10304 1372 10308
rect 1388 10364 1452 10368
rect 1388 10308 1392 10364
rect 1392 10308 1448 10364
rect 1448 10308 1452 10364
rect 1388 10304 1452 10308
rect 98932 10364 98996 10368
rect 98932 10308 98936 10364
rect 98936 10308 98992 10364
rect 98992 10308 98996 10364
rect 98932 10304 98996 10308
rect 99012 10364 99076 10368
rect 99012 10308 99016 10364
rect 99016 10308 99072 10364
rect 99072 10308 99076 10364
rect 99012 10304 99076 10308
rect 99092 10364 99156 10368
rect 99092 10308 99096 10364
rect 99096 10308 99152 10364
rect 99152 10308 99156 10364
rect 99092 10304 99156 10308
rect 99172 10364 99236 10368
rect 99172 10308 99176 10364
rect 99176 10308 99232 10364
rect 99232 10308 99236 10364
rect 99172 10304 99236 10308
rect 1676 9820 1740 9824
rect 1676 9764 1680 9820
rect 1680 9764 1736 9820
rect 1736 9764 1740 9820
rect 1676 9760 1740 9764
rect 1756 9820 1820 9824
rect 1756 9764 1760 9820
rect 1760 9764 1816 9820
rect 1816 9764 1820 9820
rect 1756 9760 1820 9764
rect 99668 9820 99732 9824
rect 99668 9764 99672 9820
rect 99672 9764 99728 9820
rect 99728 9764 99732 9820
rect 99668 9760 99732 9764
rect 99748 9820 99812 9824
rect 99748 9764 99752 9820
rect 99752 9764 99808 9820
rect 99808 9764 99812 9820
rect 99748 9760 99812 9764
rect 99828 9820 99892 9824
rect 99828 9764 99832 9820
rect 99832 9764 99888 9820
rect 99888 9764 99892 9820
rect 99828 9760 99892 9764
rect 99908 9820 99972 9824
rect 99908 9764 99912 9820
rect 99912 9764 99968 9820
rect 99968 9764 99972 9820
rect 99908 9760 99972 9764
rect 1308 9276 1372 9280
rect 1308 9220 1312 9276
rect 1312 9220 1368 9276
rect 1368 9220 1372 9276
rect 1308 9216 1372 9220
rect 1388 9276 1452 9280
rect 1388 9220 1392 9276
rect 1392 9220 1448 9276
rect 1448 9220 1452 9276
rect 1388 9216 1452 9220
rect 98932 9276 98996 9280
rect 98932 9220 98936 9276
rect 98936 9220 98992 9276
rect 98992 9220 98996 9276
rect 98932 9216 98996 9220
rect 99012 9276 99076 9280
rect 99012 9220 99016 9276
rect 99016 9220 99072 9276
rect 99072 9220 99076 9276
rect 99012 9216 99076 9220
rect 99092 9276 99156 9280
rect 99092 9220 99096 9276
rect 99096 9220 99152 9276
rect 99152 9220 99156 9276
rect 99092 9216 99156 9220
rect 99172 9276 99236 9280
rect 99172 9220 99176 9276
rect 99176 9220 99232 9276
rect 99232 9220 99236 9276
rect 99172 9216 99236 9220
rect 1676 8732 1740 8736
rect 1676 8676 1680 8732
rect 1680 8676 1736 8732
rect 1736 8676 1740 8732
rect 1676 8672 1740 8676
rect 1756 8732 1820 8736
rect 1756 8676 1760 8732
rect 1760 8676 1816 8732
rect 1816 8676 1820 8732
rect 1756 8672 1820 8676
rect 99668 8732 99732 8736
rect 99668 8676 99672 8732
rect 99672 8676 99728 8732
rect 99728 8676 99732 8732
rect 99668 8672 99732 8676
rect 99748 8732 99812 8736
rect 99748 8676 99752 8732
rect 99752 8676 99808 8732
rect 99808 8676 99812 8732
rect 99748 8672 99812 8676
rect 99828 8732 99892 8736
rect 99828 8676 99832 8732
rect 99832 8676 99888 8732
rect 99888 8676 99892 8732
rect 99828 8672 99892 8676
rect 99908 8732 99972 8736
rect 99908 8676 99912 8732
rect 99912 8676 99968 8732
rect 99968 8676 99972 8732
rect 99908 8672 99972 8676
rect 1308 8188 1372 8192
rect 1308 8132 1312 8188
rect 1312 8132 1368 8188
rect 1368 8132 1372 8188
rect 1308 8128 1372 8132
rect 1388 8188 1452 8192
rect 1388 8132 1392 8188
rect 1392 8132 1448 8188
rect 1448 8132 1452 8188
rect 1388 8128 1452 8132
rect 98932 8188 98996 8192
rect 98932 8132 98936 8188
rect 98936 8132 98992 8188
rect 98992 8132 98996 8188
rect 98932 8128 98996 8132
rect 99012 8188 99076 8192
rect 99012 8132 99016 8188
rect 99016 8132 99072 8188
rect 99072 8132 99076 8188
rect 99012 8128 99076 8132
rect 99092 8188 99156 8192
rect 99092 8132 99096 8188
rect 99096 8132 99152 8188
rect 99152 8132 99156 8188
rect 99092 8128 99156 8132
rect 99172 8188 99236 8192
rect 99172 8132 99176 8188
rect 99176 8132 99232 8188
rect 99232 8132 99236 8188
rect 99172 8128 99236 8132
rect 1676 7644 1740 7648
rect 1676 7588 1680 7644
rect 1680 7588 1736 7644
rect 1736 7588 1740 7644
rect 1676 7584 1740 7588
rect 1756 7644 1820 7648
rect 1756 7588 1760 7644
rect 1760 7588 1816 7644
rect 1816 7588 1820 7644
rect 1756 7584 1820 7588
rect 99668 7644 99732 7648
rect 99668 7588 99672 7644
rect 99672 7588 99728 7644
rect 99728 7588 99732 7644
rect 99668 7584 99732 7588
rect 99748 7644 99812 7648
rect 99748 7588 99752 7644
rect 99752 7588 99808 7644
rect 99808 7588 99812 7644
rect 99748 7584 99812 7588
rect 99828 7644 99892 7648
rect 99828 7588 99832 7644
rect 99832 7588 99888 7644
rect 99888 7588 99892 7644
rect 99828 7584 99892 7588
rect 99908 7644 99972 7648
rect 99908 7588 99912 7644
rect 99912 7588 99968 7644
rect 99968 7588 99972 7644
rect 99908 7584 99972 7588
rect 1308 7100 1372 7104
rect 1308 7044 1312 7100
rect 1312 7044 1368 7100
rect 1368 7044 1372 7100
rect 1308 7040 1372 7044
rect 1388 7100 1452 7104
rect 1388 7044 1392 7100
rect 1392 7044 1448 7100
rect 1448 7044 1452 7100
rect 1388 7040 1452 7044
rect 98932 7100 98996 7104
rect 98932 7044 98936 7100
rect 98936 7044 98992 7100
rect 98992 7044 98996 7100
rect 98932 7040 98996 7044
rect 99012 7100 99076 7104
rect 99012 7044 99016 7100
rect 99016 7044 99072 7100
rect 99072 7044 99076 7100
rect 99012 7040 99076 7044
rect 99092 7100 99156 7104
rect 99092 7044 99096 7100
rect 99096 7044 99152 7100
rect 99152 7044 99156 7100
rect 99092 7040 99156 7044
rect 99172 7100 99236 7104
rect 99172 7044 99176 7100
rect 99176 7044 99232 7100
rect 99232 7044 99236 7100
rect 99172 7040 99236 7044
rect 1676 6556 1740 6560
rect 1676 6500 1680 6556
rect 1680 6500 1736 6556
rect 1736 6500 1740 6556
rect 1676 6496 1740 6500
rect 1756 6556 1820 6560
rect 1756 6500 1760 6556
rect 1760 6500 1816 6556
rect 1816 6500 1820 6556
rect 1756 6496 1820 6500
rect 99668 6556 99732 6560
rect 99668 6500 99672 6556
rect 99672 6500 99728 6556
rect 99728 6500 99732 6556
rect 99668 6496 99732 6500
rect 99748 6556 99812 6560
rect 99748 6500 99752 6556
rect 99752 6500 99808 6556
rect 99808 6500 99812 6556
rect 99748 6496 99812 6500
rect 99828 6556 99892 6560
rect 99828 6500 99832 6556
rect 99832 6500 99888 6556
rect 99888 6500 99892 6556
rect 99828 6496 99892 6500
rect 99908 6556 99972 6560
rect 99908 6500 99912 6556
rect 99912 6500 99968 6556
rect 99968 6500 99972 6556
rect 99908 6496 99972 6500
rect 1308 6012 1372 6016
rect 1308 5956 1312 6012
rect 1312 5956 1368 6012
rect 1368 5956 1372 6012
rect 1308 5952 1372 5956
rect 1388 6012 1452 6016
rect 1388 5956 1392 6012
rect 1392 5956 1448 6012
rect 1448 5956 1452 6012
rect 1388 5952 1452 5956
rect 98932 6012 98996 6016
rect 98932 5956 98936 6012
rect 98936 5956 98992 6012
rect 98992 5956 98996 6012
rect 98932 5952 98996 5956
rect 99012 6012 99076 6016
rect 99012 5956 99016 6012
rect 99016 5956 99072 6012
rect 99072 5956 99076 6012
rect 99012 5952 99076 5956
rect 99092 6012 99156 6016
rect 99092 5956 99096 6012
rect 99096 5956 99152 6012
rect 99152 5956 99156 6012
rect 99092 5952 99156 5956
rect 99172 6012 99236 6016
rect 99172 5956 99176 6012
rect 99176 5956 99232 6012
rect 99232 5956 99236 6012
rect 99172 5952 99236 5956
rect 1676 5468 1740 5472
rect 1676 5412 1680 5468
rect 1680 5412 1736 5468
rect 1736 5412 1740 5468
rect 1676 5408 1740 5412
rect 1756 5468 1820 5472
rect 1756 5412 1760 5468
rect 1760 5412 1816 5468
rect 1816 5412 1820 5468
rect 1756 5408 1820 5412
rect 99668 5468 99732 5472
rect 99668 5412 99672 5468
rect 99672 5412 99728 5468
rect 99728 5412 99732 5468
rect 99668 5408 99732 5412
rect 99748 5468 99812 5472
rect 99748 5412 99752 5468
rect 99752 5412 99808 5468
rect 99808 5412 99812 5468
rect 99748 5408 99812 5412
rect 99828 5468 99892 5472
rect 99828 5412 99832 5468
rect 99832 5412 99888 5468
rect 99888 5412 99892 5468
rect 99828 5408 99892 5412
rect 99908 5468 99972 5472
rect 99908 5412 99912 5468
rect 99912 5412 99968 5468
rect 99968 5412 99972 5468
rect 99908 5408 99972 5412
rect 1308 4924 1372 4928
rect 1308 4868 1312 4924
rect 1312 4868 1368 4924
rect 1368 4868 1372 4924
rect 1308 4864 1372 4868
rect 1388 4924 1452 4928
rect 1388 4868 1392 4924
rect 1392 4868 1448 4924
rect 1448 4868 1452 4924
rect 1388 4864 1452 4868
rect 98932 4924 98996 4928
rect 98932 4868 98936 4924
rect 98936 4868 98992 4924
rect 98992 4868 98996 4924
rect 98932 4864 98996 4868
rect 99012 4924 99076 4928
rect 99012 4868 99016 4924
rect 99016 4868 99072 4924
rect 99072 4868 99076 4924
rect 99012 4864 99076 4868
rect 99092 4924 99156 4928
rect 99092 4868 99096 4924
rect 99096 4868 99152 4924
rect 99152 4868 99156 4924
rect 99092 4864 99156 4868
rect 99172 4924 99236 4928
rect 99172 4868 99176 4924
rect 99176 4868 99232 4924
rect 99232 4868 99236 4924
rect 99172 4864 99236 4868
rect 1676 4380 1740 4384
rect 1676 4324 1680 4380
rect 1680 4324 1736 4380
rect 1736 4324 1740 4380
rect 1676 4320 1740 4324
rect 1756 4380 1820 4384
rect 1756 4324 1760 4380
rect 1760 4324 1816 4380
rect 1816 4324 1820 4380
rect 1756 4320 1820 4324
rect 99668 4380 99732 4384
rect 99668 4324 99672 4380
rect 99672 4324 99728 4380
rect 99728 4324 99732 4380
rect 99668 4320 99732 4324
rect 99748 4380 99812 4384
rect 99748 4324 99752 4380
rect 99752 4324 99808 4380
rect 99808 4324 99812 4380
rect 99748 4320 99812 4324
rect 99828 4380 99892 4384
rect 99828 4324 99832 4380
rect 99832 4324 99888 4380
rect 99888 4324 99892 4380
rect 99828 4320 99892 4324
rect 99908 4380 99972 4384
rect 99908 4324 99912 4380
rect 99912 4324 99968 4380
rect 99968 4324 99972 4380
rect 99908 4320 99972 4324
rect 10058 3844 10122 3908
rect 84814 3844 84878 3908
rect 1308 3836 1372 3840
rect 1308 3780 1312 3836
rect 1312 3780 1368 3836
rect 1368 3780 1372 3836
rect 1308 3776 1372 3780
rect 1388 3836 1452 3840
rect 1388 3780 1392 3836
rect 1392 3780 1448 3836
rect 1448 3780 1452 3836
rect 1388 3776 1452 3780
rect 98932 3836 98996 3840
rect 98932 3780 98936 3836
rect 98936 3780 98992 3836
rect 98992 3780 98996 3836
rect 98932 3776 98996 3780
rect 99012 3836 99076 3840
rect 99012 3780 99016 3836
rect 99016 3780 99072 3836
rect 99072 3780 99076 3836
rect 99012 3776 99076 3780
rect 99092 3836 99156 3840
rect 99092 3780 99096 3836
rect 99096 3780 99152 3836
rect 99152 3780 99156 3836
rect 99092 3776 99156 3780
rect 99172 3836 99236 3840
rect 99172 3780 99176 3836
rect 99176 3780 99232 3836
rect 99232 3780 99236 3836
rect 99172 3776 99236 3780
rect 84665 3708 84729 3772
rect 84527 3572 84591 3636
rect 17438 3496 17502 3500
rect 17438 3440 17462 3496
rect 17462 3440 17502 3496
rect 17438 3436 17502 3440
rect 19774 3436 19838 3500
rect 20942 3436 21006 3500
rect 22110 3436 22174 3500
rect 24446 3496 24510 3500
rect 24446 3440 24490 3496
rect 24490 3440 24510 3496
rect 24446 3436 24510 3440
rect 25614 3436 25678 3500
rect 26782 3436 26846 3500
rect 27936 3436 28000 3500
rect 30286 3496 30350 3500
rect 30286 3440 30342 3496
rect 30342 3440 30350 3496
rect 30286 3436 30350 3440
rect 33790 3436 33854 3500
rect 34958 3436 35022 3500
rect 1676 3292 1740 3296
rect 1676 3236 1680 3292
rect 1680 3236 1736 3292
rect 1736 3236 1740 3292
rect 1676 3232 1740 3236
rect 1756 3292 1820 3296
rect 1756 3236 1760 3292
rect 1760 3236 1816 3292
rect 1816 3236 1820 3292
rect 1756 3232 1820 3236
rect 99668 3292 99732 3296
rect 99668 3236 99672 3292
rect 99672 3236 99728 3292
rect 99728 3236 99732 3292
rect 99668 3232 99732 3236
rect 99748 3292 99812 3296
rect 99748 3236 99752 3292
rect 99752 3236 99808 3292
rect 99808 3236 99812 3292
rect 99748 3232 99812 3236
rect 99828 3292 99892 3296
rect 99828 3236 99832 3292
rect 99832 3236 99888 3292
rect 99888 3236 99892 3292
rect 99828 3232 99892 3236
rect 99908 3292 99972 3296
rect 99908 3236 99912 3292
rect 99912 3236 99968 3292
rect 99968 3236 99972 3292
rect 99908 3232 99972 3236
rect 18644 2816 18708 2820
rect 18644 2760 18694 2816
rect 18694 2760 18708 2816
rect 18644 2756 18708 2760
rect 23244 2816 23308 2820
rect 23244 2760 23258 2816
rect 23258 2760 23308 2816
rect 23244 2756 23308 2760
rect 29132 2756 29196 2820
rect 31524 2816 31588 2820
rect 31524 2760 31574 2816
rect 31574 2760 31588 2816
rect 31524 2756 31588 2760
rect 32628 2756 32692 2820
rect 36124 2816 36188 2820
rect 36124 2760 36138 2816
rect 36138 2760 36188 2816
rect 36124 2756 36188 2760
rect 37228 2756 37292 2820
rect 1308 2748 1372 2752
rect 1308 2692 1312 2748
rect 1312 2692 1368 2748
rect 1368 2692 1372 2748
rect 1308 2688 1372 2692
rect 1388 2748 1452 2752
rect 1388 2692 1392 2748
rect 1392 2692 1448 2748
rect 1448 2692 1452 2748
rect 1388 2688 1452 2692
rect 98932 2748 98996 2752
rect 98932 2692 98936 2748
rect 98936 2692 98992 2748
rect 98992 2692 98996 2748
rect 98932 2688 98996 2692
rect 99012 2748 99076 2752
rect 99012 2692 99016 2748
rect 99016 2692 99072 2748
rect 99072 2692 99076 2748
rect 99012 2688 99076 2692
rect 99092 2748 99156 2752
rect 99092 2692 99096 2748
rect 99096 2692 99152 2748
rect 99152 2692 99156 2748
rect 99092 2688 99156 2692
rect 99172 2748 99236 2752
rect 99172 2692 99176 2748
rect 99176 2692 99232 2748
rect 99232 2692 99236 2748
rect 99172 2688 99236 2692
rect 1676 2204 1740 2208
rect 1676 2148 1680 2204
rect 1680 2148 1736 2204
rect 1736 2148 1740 2204
rect 1676 2144 1740 2148
rect 1756 2204 1820 2208
rect 1756 2148 1760 2204
rect 1760 2148 1816 2204
rect 1816 2148 1820 2204
rect 1756 2144 1820 2148
rect 99668 2204 99732 2208
rect 99668 2148 99672 2204
rect 99672 2148 99728 2204
rect 99728 2148 99732 2204
rect 99668 2144 99732 2148
rect 99748 2204 99812 2208
rect 99748 2148 99752 2204
rect 99752 2148 99808 2204
rect 99808 2148 99812 2204
rect 99748 2144 99812 2148
rect 99828 2204 99892 2208
rect 99828 2148 99832 2204
rect 99832 2148 99888 2204
rect 99888 2148 99892 2204
rect 99828 2144 99892 2148
rect 99908 2204 99972 2208
rect 99908 2148 99912 2204
rect 99912 2148 99968 2204
rect 99968 2148 99972 2204
rect 99908 2144 99972 2148
<< metal4 >>
rect 4208 101760 4528 101776
rect 4208 101696 4216 101760
rect 4280 101696 4296 101760
rect 4360 101696 4376 101760
rect 4440 101696 4456 101760
rect 4520 101696 4528 101760
rect 4208 100672 4528 101696
rect 4208 100608 4216 100672
rect 4280 100608 4296 100672
rect 4360 100608 4376 100672
rect 4440 100608 4456 100672
rect 4520 100608 4528 100672
rect 4208 99584 4528 100608
rect 4208 99520 4216 99584
rect 4280 99520 4296 99584
rect 4360 99520 4376 99584
rect 4440 99520 4456 99584
rect 4520 99520 4528 99584
rect 4208 98496 4528 99520
rect 4208 98432 4216 98496
rect 4280 98432 4296 98496
rect 4360 98432 4376 98496
rect 4440 98432 4456 98496
rect 4520 98432 4528 98496
rect 4208 97532 4528 98432
rect 4208 97408 4250 97532
rect 4486 97408 4528 97532
rect 4208 97344 4216 97408
rect 4520 97344 4528 97408
rect 4208 97296 4250 97344
rect 4486 97296 4528 97344
rect 4208 96320 4528 97296
rect 4208 96256 4216 96320
rect 4280 96256 4296 96320
rect 4360 96256 4376 96320
rect 4440 96256 4456 96320
rect 4520 96256 4528 96320
rect 4208 95232 4528 96256
rect 4208 95168 4216 95232
rect 4280 95168 4296 95232
rect 4360 95168 4376 95232
rect 4440 95168 4456 95232
rect 4520 95168 4528 95232
rect 4208 94144 4528 95168
rect 4208 94080 4216 94144
rect 4280 94080 4296 94144
rect 4360 94080 4376 94144
rect 4440 94080 4456 94144
rect 4520 94080 4528 94144
rect 4208 93056 4528 94080
rect 4208 92992 4216 93056
rect 4280 92992 4296 93056
rect 4360 92992 4376 93056
rect 4440 92992 4456 93056
rect 4520 92992 4528 93056
rect 4208 91968 4528 92992
rect 4208 91904 4216 91968
rect 4280 91904 4296 91968
rect 4360 91904 4376 91968
rect 4440 91904 4456 91968
rect 4520 91904 4528 91968
rect 4208 90880 4528 91904
rect 4208 90816 4216 90880
rect 4280 90816 4296 90880
rect 4360 90816 4376 90880
rect 4440 90816 4456 90880
rect 4520 90816 4528 90880
rect 4208 89792 4528 90816
rect 4208 89728 4216 89792
rect 4280 89728 4296 89792
rect 4360 89728 4376 89792
rect 4440 89728 4456 89792
rect 4520 89728 4528 89792
rect 4208 88704 4528 89728
rect 4208 88640 4216 88704
rect 4280 88640 4296 88704
rect 4360 88640 4376 88704
rect 4440 88640 4456 88704
rect 4520 88640 4528 88704
rect 4208 87616 4528 88640
rect 4208 87552 4216 87616
rect 4280 87552 4296 87616
rect 4360 87552 4376 87616
rect 4440 87552 4456 87616
rect 4520 87552 4528 87616
rect 4208 86528 4528 87552
rect 4208 86464 4216 86528
rect 4280 86464 4296 86528
rect 4360 86464 4376 86528
rect 4440 86464 4456 86528
rect 4520 86464 4528 86528
rect 4208 85440 4528 86464
rect 4208 85376 4216 85440
rect 4280 85376 4296 85440
rect 4360 85376 4376 85440
rect 4440 85376 4456 85440
rect 4520 85376 4528 85440
rect 4208 84352 4528 85376
rect 4208 84288 4216 84352
rect 4280 84288 4296 84352
rect 4360 84288 4376 84352
rect 4440 84288 4456 84352
rect 4520 84288 4528 84352
rect 4208 83264 4528 84288
rect 4208 83200 4216 83264
rect 4280 83200 4296 83264
rect 4360 83200 4376 83264
rect 4440 83200 4456 83264
rect 4520 83200 4528 83264
rect 4208 82176 4528 83200
rect 4208 82112 4216 82176
rect 4280 82112 4296 82176
rect 4360 82112 4376 82176
rect 4440 82112 4456 82176
rect 4520 82112 4528 82176
rect 4208 81088 4528 82112
rect 4208 81024 4216 81088
rect 4280 81024 4296 81088
rect 4360 81024 4376 81088
rect 4440 81024 4456 81088
rect 4520 81024 4528 81088
rect 4208 80000 4528 81024
rect 4208 79936 4216 80000
rect 4280 79936 4296 80000
rect 4360 79936 4376 80000
rect 4440 79936 4456 80000
rect 4520 79936 4528 80000
rect 4208 78912 4528 79936
rect 4208 78848 4216 78912
rect 4280 78848 4296 78912
rect 4360 78848 4376 78912
rect 4440 78848 4456 78912
rect 4520 78848 4528 78912
rect 4208 77824 4528 78848
rect 4208 77760 4216 77824
rect 4280 77760 4296 77824
rect 4360 77760 4376 77824
rect 4440 77760 4456 77824
rect 4520 77760 4528 77824
rect 4208 76736 4528 77760
rect 4208 76672 4216 76736
rect 4280 76672 4296 76736
rect 4360 76672 4376 76736
rect 4440 76672 4456 76736
rect 4520 76672 4528 76736
rect 4208 75648 4528 76672
rect 4208 75584 4216 75648
rect 4280 75584 4296 75648
rect 4360 75584 4376 75648
rect 4440 75584 4456 75648
rect 4520 75584 4528 75648
rect 4208 74560 4528 75584
rect 4208 74496 4216 74560
rect 4280 74496 4296 74560
rect 4360 74496 4376 74560
rect 4440 74496 4456 74560
rect 4520 74496 4528 74560
rect 4208 73472 4528 74496
rect 4208 73408 4216 73472
rect 4280 73408 4296 73472
rect 4360 73408 4376 73472
rect 4440 73408 4456 73472
rect 4520 73408 4528 73472
rect 4208 72384 4528 73408
rect 4208 72320 4216 72384
rect 4280 72320 4296 72384
rect 4360 72320 4376 72384
rect 4440 72320 4456 72384
rect 4520 72320 4528 72384
rect 4208 71296 4528 72320
rect 4208 71232 4216 71296
rect 4280 71232 4296 71296
rect 4360 71232 4376 71296
rect 4440 71232 4456 71296
rect 4520 71232 4528 71296
rect 4208 70208 4528 71232
rect 4208 70144 4216 70208
rect 4280 70144 4296 70208
rect 4360 70144 4376 70208
rect 4440 70144 4456 70208
rect 4520 70144 4528 70208
rect 4208 69120 4528 70144
rect 4208 69056 4216 69120
rect 4280 69056 4296 69120
rect 4360 69056 4376 69120
rect 4440 69056 4456 69120
rect 4520 69056 4528 69120
rect 4208 68032 4528 69056
rect 4208 67968 4216 68032
rect 4280 67968 4296 68032
rect 4360 67968 4376 68032
rect 4440 67968 4456 68032
rect 4520 67968 4528 68032
rect 4208 66944 4528 67968
rect 4208 66880 4216 66944
rect 4280 66896 4296 66944
rect 4360 66896 4376 66944
rect 4440 66896 4456 66944
rect 4520 66880 4528 66944
rect 4208 66660 4250 66880
rect 4486 66660 4528 66880
rect 4208 65856 4528 66660
rect 4208 65792 4216 65856
rect 4280 65792 4296 65856
rect 4360 65792 4376 65856
rect 4440 65792 4456 65856
rect 4520 65792 4528 65856
rect 4208 64768 4528 65792
rect 4208 64704 4216 64768
rect 4280 64704 4296 64768
rect 4360 64704 4376 64768
rect 4440 64704 4456 64768
rect 4520 64704 4528 64768
rect 4208 63680 4528 64704
rect 4208 63616 4216 63680
rect 4280 63616 4296 63680
rect 4360 63616 4376 63680
rect 4440 63616 4456 63680
rect 4520 63616 4528 63680
rect 4208 62592 4528 63616
rect 4208 62528 4216 62592
rect 4280 62528 4296 62592
rect 4360 62528 4376 62592
rect 4440 62528 4456 62592
rect 4520 62528 4528 62592
rect 4208 61504 4528 62528
rect 4208 61440 4216 61504
rect 4280 61440 4296 61504
rect 4360 61440 4376 61504
rect 4440 61440 4456 61504
rect 4520 61440 4528 61504
rect 1300 60416 1460 60432
rect 1300 60352 1308 60416
rect 1372 60352 1388 60416
rect 1452 60352 1460 60416
rect 1300 59328 1460 60352
rect 1300 59264 1308 59328
rect 1372 59264 1388 59328
rect 1452 59264 1460 59328
rect 1300 58240 1460 59264
rect 1300 58176 1308 58240
rect 1372 58176 1388 58240
rect 1452 58176 1460 58240
rect 1300 57152 1460 58176
rect 1300 57088 1308 57152
rect 1372 57088 1388 57152
rect 1452 57088 1460 57152
rect 1300 56064 1460 57088
rect 1300 56000 1308 56064
rect 1372 56000 1388 56064
rect 1452 56000 1460 56064
rect 1300 54976 1460 56000
rect 1300 54912 1308 54976
rect 1372 54912 1388 54976
rect 1452 54912 1460 54976
rect 1300 53888 1460 54912
rect 1300 53824 1308 53888
rect 1372 53824 1388 53888
rect 1452 53824 1460 53888
rect 1300 52800 1460 53824
rect 1300 52736 1308 52800
rect 1372 52736 1388 52800
rect 1452 52736 1460 52800
rect 1300 51712 1460 52736
rect 1300 51648 1308 51712
rect 1372 51648 1388 51712
rect 1452 51648 1460 51712
rect 1300 50624 1460 51648
rect 1300 50560 1308 50624
rect 1372 50560 1388 50624
rect 1452 50560 1460 50624
rect 1300 49536 1460 50560
rect 1300 49472 1308 49536
rect 1372 49472 1388 49536
rect 1452 49472 1460 49536
rect 1300 48448 1460 49472
rect 1300 48384 1308 48448
rect 1372 48384 1388 48448
rect 1452 48384 1460 48448
rect 1300 47360 1460 48384
rect 1300 47296 1308 47360
rect 1372 47296 1388 47360
rect 1452 47296 1460 47360
rect 1300 46272 1460 47296
rect 1300 46208 1308 46272
rect 1372 46208 1388 46272
rect 1452 46208 1460 46272
rect 1300 45184 1460 46208
rect 1300 45120 1308 45184
rect 1372 45120 1388 45184
rect 1452 45120 1460 45184
rect 1300 44096 1460 45120
rect 1300 44032 1308 44096
rect 1372 44032 1388 44096
rect 1452 44032 1460 44096
rect 1300 43008 1460 44032
rect 1300 42944 1308 43008
rect 1372 42944 1388 43008
rect 1452 42944 1460 43008
rect 1300 41920 1460 42944
rect 1300 41856 1308 41920
rect 1372 41856 1388 41920
rect 1452 41856 1460 41920
rect 1300 40832 1460 41856
rect 1300 40768 1308 40832
rect 1372 40768 1388 40832
rect 1452 40768 1460 40832
rect 1300 39744 1460 40768
rect 1300 39680 1308 39744
rect 1372 39680 1388 39744
rect 1452 39680 1460 39744
rect 1300 38656 1460 39680
rect 1300 38592 1308 38656
rect 1372 38592 1388 38656
rect 1452 38592 1460 38656
rect 1300 37568 1460 38592
rect 1300 37504 1308 37568
rect 1372 37504 1388 37568
rect 1452 37504 1460 37568
rect 1300 36480 1460 37504
rect 1300 36416 1308 36480
rect 1372 36416 1388 36480
rect 1452 36416 1460 36480
rect 1300 35392 1460 36416
rect 1300 35328 1308 35392
rect 1372 35328 1388 35392
rect 1452 35328 1460 35392
rect 1300 34304 1460 35328
rect 1300 34240 1308 34304
rect 1372 34240 1388 34304
rect 1452 34240 1460 34304
rect 1300 33216 1460 34240
rect 1300 33152 1308 33216
rect 1372 33152 1388 33216
rect 1452 33152 1460 33216
rect 1300 32128 1460 33152
rect 1300 32064 1308 32128
rect 1372 32064 1388 32128
rect 1452 32064 1460 32128
rect 1300 31040 1460 32064
rect 1300 30976 1308 31040
rect 1372 30976 1388 31040
rect 1452 30976 1460 31040
rect 1300 29952 1460 30976
rect 1300 29888 1308 29952
rect 1372 29888 1388 29952
rect 1452 29888 1460 29952
rect 1300 28864 1460 29888
rect 1300 28800 1308 28864
rect 1372 28800 1388 28864
rect 1452 28800 1460 28864
rect 1300 27776 1460 28800
rect 1300 27712 1308 27776
rect 1372 27712 1388 27776
rect 1452 27712 1460 27776
rect 1300 26688 1460 27712
rect 1300 26624 1308 26688
rect 1372 26624 1388 26688
rect 1452 26624 1460 26688
rect 1300 25600 1460 26624
rect 1300 25536 1308 25600
rect 1372 25536 1388 25600
rect 1452 25536 1460 25600
rect 1300 24512 1460 25536
rect 1300 24448 1308 24512
rect 1372 24448 1388 24512
rect 1452 24448 1460 24512
rect 1300 23424 1460 24448
rect 1300 23360 1308 23424
rect 1372 23360 1388 23424
rect 1452 23360 1460 23424
rect 1300 22336 1460 23360
rect 1300 22272 1308 22336
rect 1372 22272 1388 22336
rect 1452 22272 1460 22336
rect 1300 21248 1460 22272
rect 1300 21184 1308 21248
rect 1372 21184 1388 21248
rect 1452 21184 1460 21248
rect 1300 20160 1460 21184
rect 1300 20096 1308 20160
rect 1372 20096 1388 20160
rect 1452 20096 1460 20160
rect 1300 19072 1460 20096
rect 1300 19008 1308 19072
rect 1372 19008 1388 19072
rect 1452 19008 1460 19072
rect 1300 17984 1460 19008
rect 1300 17920 1308 17984
rect 1372 17920 1388 17984
rect 1452 17920 1460 17984
rect 1300 16896 1460 17920
rect 1300 16832 1308 16896
rect 1372 16832 1388 16896
rect 1452 16832 1460 16896
rect 1300 15808 1460 16832
rect 1300 15744 1308 15808
rect 1372 15744 1388 15808
rect 1452 15744 1460 15808
rect 1300 14720 1460 15744
rect 1300 14656 1308 14720
rect 1372 14656 1388 14720
rect 1452 14656 1460 14720
rect 1300 13632 1460 14656
rect 1300 13568 1308 13632
rect 1372 13568 1388 13632
rect 1452 13568 1460 13632
rect 1300 12544 1460 13568
rect 1300 12480 1308 12544
rect 1372 12480 1388 12544
rect 1452 12480 1460 12544
rect 1300 11456 1460 12480
rect 1300 11392 1308 11456
rect 1372 11392 1388 11456
rect 1452 11392 1460 11456
rect 1300 10368 1460 11392
rect 1300 10304 1308 10368
rect 1372 10304 1388 10368
rect 1452 10304 1460 10368
rect 1300 9280 1460 10304
rect 1300 9216 1308 9280
rect 1372 9216 1388 9280
rect 1452 9216 1460 9280
rect 1300 8192 1460 9216
rect 1300 8128 1308 8192
rect 1372 8128 1388 8192
rect 1452 8128 1460 8192
rect 1300 7104 1460 8128
rect 1300 7040 1308 7104
rect 1372 7040 1388 7104
rect 1452 7040 1460 7104
rect 1300 6016 1460 7040
rect 1300 5952 1308 6016
rect 1372 5952 1388 6016
rect 1452 5952 1460 6016
rect 1300 4928 1460 5952
rect 1300 4864 1308 4928
rect 1372 4864 1388 4928
rect 1452 4864 1460 4928
rect 1300 3840 1460 4864
rect 1300 3776 1308 3840
rect 1372 3776 1388 3840
rect 1452 3776 1460 3840
rect 1300 2752 1460 3776
rect 1300 2688 1308 2752
rect 1372 2688 1388 2752
rect 1452 2688 1460 2752
rect 1300 2128 1460 2688
rect 1668 59872 1828 60432
rect 1668 59808 1676 59872
rect 1740 59808 1756 59872
rect 1820 59808 1828 59872
rect 4208 60416 4528 61440
rect 4208 60352 4216 60416
rect 4280 60352 4296 60416
rect 4360 60352 4376 60416
rect 4440 60352 4456 60416
rect 4520 60352 4528 60416
rect 4208 59834 4528 60352
rect 4868 101216 5188 101776
rect 4868 101152 4876 101216
rect 4940 101152 4956 101216
rect 5020 101152 5036 101216
rect 5100 101152 5116 101216
rect 5180 101152 5188 101216
rect 4868 100128 5188 101152
rect 4868 100064 4876 100128
rect 4940 100064 4956 100128
rect 5020 100064 5036 100128
rect 5100 100064 5116 100128
rect 5180 100064 5188 100128
rect 4868 99040 5188 100064
rect 4868 98976 4876 99040
rect 4940 98976 4956 99040
rect 5020 98976 5036 99040
rect 5100 98976 5116 99040
rect 5180 98976 5188 99040
rect 4868 98192 5188 98976
rect 4868 97956 4910 98192
rect 5146 97956 5188 98192
rect 4868 97952 5188 97956
rect 4868 97888 4876 97952
rect 4940 97888 4956 97952
rect 5020 97888 5036 97952
rect 5100 97888 5116 97952
rect 5180 97888 5188 97952
rect 4868 96864 5188 97888
rect 4868 96800 4876 96864
rect 4940 96800 4956 96864
rect 5020 96800 5036 96864
rect 5100 96800 5116 96864
rect 5180 96800 5188 96864
rect 4868 95776 5188 96800
rect 4868 95712 4876 95776
rect 4940 95712 4956 95776
rect 5020 95712 5036 95776
rect 5100 95712 5116 95776
rect 5180 95712 5188 95776
rect 4868 94688 5188 95712
rect 4868 94624 4876 94688
rect 4940 94624 4956 94688
rect 5020 94624 5036 94688
rect 5100 94624 5116 94688
rect 5180 94624 5188 94688
rect 4868 93600 5188 94624
rect 4868 93536 4876 93600
rect 4940 93536 4956 93600
rect 5020 93536 5036 93600
rect 5100 93536 5116 93600
rect 5180 93536 5188 93600
rect 4868 92512 5188 93536
rect 4868 92448 4876 92512
rect 4940 92448 4956 92512
rect 5020 92448 5036 92512
rect 5100 92448 5116 92512
rect 5180 92448 5188 92512
rect 4868 91424 5188 92448
rect 4868 91360 4876 91424
rect 4940 91360 4956 91424
rect 5020 91360 5036 91424
rect 5100 91360 5116 91424
rect 5180 91360 5188 91424
rect 4868 90336 5188 91360
rect 4868 90272 4876 90336
rect 4940 90272 4956 90336
rect 5020 90272 5036 90336
rect 5100 90272 5116 90336
rect 5180 90272 5188 90336
rect 4868 89248 5188 90272
rect 4868 89184 4876 89248
rect 4940 89184 4956 89248
rect 5020 89184 5036 89248
rect 5100 89184 5116 89248
rect 5180 89184 5188 89248
rect 4868 88160 5188 89184
rect 4868 88096 4876 88160
rect 4940 88096 4956 88160
rect 5020 88096 5036 88160
rect 5100 88096 5116 88160
rect 5180 88096 5188 88160
rect 4868 87072 5188 88096
rect 4868 87008 4876 87072
rect 4940 87008 4956 87072
rect 5020 87008 5036 87072
rect 5100 87008 5116 87072
rect 5180 87008 5188 87072
rect 4868 85984 5188 87008
rect 4868 85920 4876 85984
rect 4940 85920 4956 85984
rect 5020 85920 5036 85984
rect 5100 85920 5116 85984
rect 5180 85920 5188 85984
rect 4868 84896 5188 85920
rect 4868 84832 4876 84896
rect 4940 84832 4956 84896
rect 5020 84832 5036 84896
rect 5100 84832 5116 84896
rect 5180 84832 5188 84896
rect 4868 83808 5188 84832
rect 4868 83744 4876 83808
rect 4940 83744 4956 83808
rect 5020 83744 5036 83808
rect 5100 83744 5116 83808
rect 5180 83744 5188 83808
rect 4868 82720 5188 83744
rect 4868 82656 4876 82720
rect 4940 82656 4956 82720
rect 5020 82656 5036 82720
rect 5100 82656 5116 82720
rect 5180 82656 5188 82720
rect 4868 81632 5188 82656
rect 4868 81568 4876 81632
rect 4940 81568 4956 81632
rect 5020 81568 5036 81632
rect 5100 81568 5116 81632
rect 5180 81568 5188 81632
rect 4868 80544 5188 81568
rect 4868 80480 4876 80544
rect 4940 80480 4956 80544
rect 5020 80480 5036 80544
rect 5100 80480 5116 80544
rect 5180 80480 5188 80544
rect 4868 79456 5188 80480
rect 4868 79392 4876 79456
rect 4940 79392 4956 79456
rect 5020 79392 5036 79456
rect 5100 79392 5116 79456
rect 5180 79392 5188 79456
rect 4868 78368 5188 79392
rect 4868 78304 4876 78368
rect 4940 78304 4956 78368
rect 5020 78304 5036 78368
rect 5100 78304 5116 78368
rect 5180 78304 5188 78368
rect 4868 77280 5188 78304
rect 4868 77216 4876 77280
rect 4940 77216 4956 77280
rect 5020 77216 5036 77280
rect 5100 77216 5116 77280
rect 5180 77216 5188 77280
rect 4868 76192 5188 77216
rect 4868 76128 4876 76192
rect 4940 76128 4956 76192
rect 5020 76128 5036 76192
rect 5100 76128 5116 76192
rect 5180 76128 5188 76192
rect 4868 75104 5188 76128
rect 4868 75040 4876 75104
rect 4940 75040 4956 75104
rect 5020 75040 5036 75104
rect 5100 75040 5116 75104
rect 5180 75040 5188 75104
rect 4868 74016 5188 75040
rect 4868 73952 4876 74016
rect 4940 73952 4956 74016
rect 5020 73952 5036 74016
rect 5100 73952 5116 74016
rect 5180 73952 5188 74016
rect 4868 72928 5188 73952
rect 4868 72864 4876 72928
rect 4940 72864 4956 72928
rect 5020 72864 5036 72928
rect 5100 72864 5116 72928
rect 5180 72864 5188 72928
rect 4868 71840 5188 72864
rect 4868 71776 4876 71840
rect 4940 71776 4956 71840
rect 5020 71776 5036 71840
rect 5100 71776 5116 71840
rect 5180 71776 5188 71840
rect 4868 70752 5188 71776
rect 4868 70688 4876 70752
rect 4940 70688 4956 70752
rect 5020 70688 5036 70752
rect 5100 70688 5116 70752
rect 5180 70688 5188 70752
rect 4868 69664 5188 70688
rect 4868 69600 4876 69664
rect 4940 69600 4956 69664
rect 5020 69600 5036 69664
rect 5100 69600 5116 69664
rect 5180 69600 5188 69664
rect 4868 68576 5188 69600
rect 4868 68512 4876 68576
rect 4940 68512 4956 68576
rect 5020 68512 5036 68576
rect 5100 68512 5116 68576
rect 5180 68512 5188 68576
rect 4868 67556 5188 68512
rect 4868 67488 4910 67556
rect 5146 67488 5188 67556
rect 4868 67424 4876 67488
rect 5180 67424 5188 67488
rect 4868 67320 4910 67424
rect 5146 67320 5188 67424
rect 4868 66400 5188 67320
rect 4868 66336 4876 66400
rect 4940 66336 4956 66400
rect 5020 66336 5036 66400
rect 5100 66336 5116 66400
rect 5180 66336 5188 66400
rect 4868 65312 5188 66336
rect 4868 65248 4876 65312
rect 4940 65248 4956 65312
rect 5020 65248 5036 65312
rect 5100 65248 5116 65312
rect 5180 65248 5188 65312
rect 4868 64224 5188 65248
rect 4868 64160 4876 64224
rect 4940 64160 4956 64224
rect 5020 64160 5036 64224
rect 5100 64160 5116 64224
rect 5180 64160 5188 64224
rect 4868 63136 5188 64160
rect 4868 63072 4876 63136
rect 4940 63072 4956 63136
rect 5020 63072 5036 63136
rect 5100 63072 5116 63136
rect 5180 63072 5188 63136
rect 4868 62048 5188 63072
rect 4868 61984 4876 62048
rect 4940 61984 4956 62048
rect 5020 61984 5036 62048
rect 5100 61984 5116 62048
rect 5180 61984 5188 62048
rect 4868 60960 5188 61984
rect 4868 60896 4876 60960
rect 4940 60896 4956 60960
rect 5020 60896 5036 60960
rect 5100 60896 5116 60960
rect 5180 60896 5188 60960
rect 4868 59872 5188 60896
rect 1668 58784 1828 59808
rect 4868 59808 4876 59872
rect 4940 59808 4956 59872
rect 5020 59808 5036 59872
rect 5100 59808 5116 59872
rect 5180 59808 5188 59872
rect 34928 101760 35248 101776
rect 34928 101696 34936 101760
rect 35000 101696 35016 101760
rect 35080 101696 35096 101760
rect 35160 101696 35176 101760
rect 35240 101696 35248 101760
rect 34928 100672 35248 101696
rect 34928 100608 34936 100672
rect 35000 100608 35016 100672
rect 35080 100608 35096 100672
rect 35160 100608 35176 100672
rect 35240 100608 35248 100672
rect 34928 99584 35248 100608
rect 34928 99520 34936 99584
rect 35000 99520 35016 99584
rect 35080 99520 35096 99584
rect 35160 99520 35176 99584
rect 35240 99520 35248 99584
rect 34928 98496 35248 99520
rect 34928 98432 34936 98496
rect 35000 98432 35016 98496
rect 35080 98432 35096 98496
rect 35160 98432 35176 98496
rect 35240 98432 35248 98496
rect 34928 97532 35248 98432
rect 34928 97408 34970 97532
rect 35206 97408 35248 97532
rect 34928 97344 34936 97408
rect 35240 97344 35248 97408
rect 34928 97296 34970 97344
rect 35206 97296 35248 97344
rect 34928 96320 35248 97296
rect 34928 96256 34936 96320
rect 35000 96256 35016 96320
rect 35080 96256 35096 96320
rect 35160 96256 35176 96320
rect 35240 96256 35248 96320
rect 34928 95232 35248 96256
rect 34928 95168 34936 95232
rect 35000 95168 35016 95232
rect 35080 95168 35096 95232
rect 35160 95168 35176 95232
rect 35240 95168 35248 95232
rect 34928 94144 35248 95168
rect 34928 94080 34936 94144
rect 35000 94080 35016 94144
rect 35080 94080 35096 94144
rect 35160 94080 35176 94144
rect 35240 94080 35248 94144
rect 34928 93056 35248 94080
rect 34928 92992 34936 93056
rect 35000 92992 35016 93056
rect 35080 92992 35096 93056
rect 35160 92992 35176 93056
rect 35240 92992 35248 93056
rect 34928 91968 35248 92992
rect 34928 91904 34936 91968
rect 35000 91904 35016 91968
rect 35080 91904 35096 91968
rect 35160 91904 35176 91968
rect 35240 91904 35248 91968
rect 34928 90880 35248 91904
rect 34928 90816 34936 90880
rect 35000 90816 35016 90880
rect 35080 90816 35096 90880
rect 35160 90816 35176 90880
rect 35240 90816 35248 90880
rect 34928 89792 35248 90816
rect 34928 89728 34936 89792
rect 35000 89728 35016 89792
rect 35080 89728 35096 89792
rect 35160 89728 35176 89792
rect 35240 89728 35248 89792
rect 34928 88704 35248 89728
rect 34928 88640 34936 88704
rect 35000 88640 35016 88704
rect 35080 88640 35096 88704
rect 35160 88640 35176 88704
rect 35240 88640 35248 88704
rect 34928 87616 35248 88640
rect 34928 87552 34936 87616
rect 35000 87552 35016 87616
rect 35080 87552 35096 87616
rect 35160 87552 35176 87616
rect 35240 87552 35248 87616
rect 34928 86528 35248 87552
rect 34928 86464 34936 86528
rect 35000 86464 35016 86528
rect 35080 86464 35096 86528
rect 35160 86464 35176 86528
rect 35240 86464 35248 86528
rect 34928 85440 35248 86464
rect 34928 85376 34936 85440
rect 35000 85376 35016 85440
rect 35080 85376 35096 85440
rect 35160 85376 35176 85440
rect 35240 85376 35248 85440
rect 34928 84352 35248 85376
rect 34928 84288 34936 84352
rect 35000 84288 35016 84352
rect 35080 84288 35096 84352
rect 35160 84288 35176 84352
rect 35240 84288 35248 84352
rect 34928 83264 35248 84288
rect 34928 83200 34936 83264
rect 35000 83200 35016 83264
rect 35080 83200 35096 83264
rect 35160 83200 35176 83264
rect 35240 83200 35248 83264
rect 34928 82176 35248 83200
rect 34928 82112 34936 82176
rect 35000 82112 35016 82176
rect 35080 82112 35096 82176
rect 35160 82112 35176 82176
rect 35240 82112 35248 82176
rect 34928 81088 35248 82112
rect 34928 81024 34936 81088
rect 35000 81024 35016 81088
rect 35080 81024 35096 81088
rect 35160 81024 35176 81088
rect 35240 81024 35248 81088
rect 34928 80000 35248 81024
rect 34928 79936 34936 80000
rect 35000 79936 35016 80000
rect 35080 79936 35096 80000
rect 35160 79936 35176 80000
rect 35240 79936 35248 80000
rect 34928 78912 35248 79936
rect 34928 78848 34936 78912
rect 35000 78848 35016 78912
rect 35080 78848 35096 78912
rect 35160 78848 35176 78912
rect 35240 78848 35248 78912
rect 34928 77824 35248 78848
rect 34928 77760 34936 77824
rect 35000 77760 35016 77824
rect 35080 77760 35096 77824
rect 35160 77760 35176 77824
rect 35240 77760 35248 77824
rect 34928 76736 35248 77760
rect 34928 76672 34936 76736
rect 35000 76672 35016 76736
rect 35080 76672 35096 76736
rect 35160 76672 35176 76736
rect 35240 76672 35248 76736
rect 34928 75648 35248 76672
rect 34928 75584 34936 75648
rect 35000 75584 35016 75648
rect 35080 75584 35096 75648
rect 35160 75584 35176 75648
rect 35240 75584 35248 75648
rect 34928 74560 35248 75584
rect 34928 74496 34936 74560
rect 35000 74496 35016 74560
rect 35080 74496 35096 74560
rect 35160 74496 35176 74560
rect 35240 74496 35248 74560
rect 34928 73472 35248 74496
rect 34928 73408 34936 73472
rect 35000 73408 35016 73472
rect 35080 73408 35096 73472
rect 35160 73408 35176 73472
rect 35240 73408 35248 73472
rect 34928 72384 35248 73408
rect 34928 72320 34936 72384
rect 35000 72320 35016 72384
rect 35080 72320 35096 72384
rect 35160 72320 35176 72384
rect 35240 72320 35248 72384
rect 34928 71296 35248 72320
rect 34928 71232 34936 71296
rect 35000 71232 35016 71296
rect 35080 71232 35096 71296
rect 35160 71232 35176 71296
rect 35240 71232 35248 71296
rect 34928 70208 35248 71232
rect 34928 70144 34936 70208
rect 35000 70144 35016 70208
rect 35080 70144 35096 70208
rect 35160 70144 35176 70208
rect 35240 70144 35248 70208
rect 34928 69120 35248 70144
rect 34928 69056 34936 69120
rect 35000 69056 35016 69120
rect 35080 69056 35096 69120
rect 35160 69056 35176 69120
rect 35240 69056 35248 69120
rect 34928 68032 35248 69056
rect 34928 67968 34936 68032
rect 35000 67968 35016 68032
rect 35080 67968 35096 68032
rect 35160 67968 35176 68032
rect 35240 67968 35248 68032
rect 34928 66944 35248 67968
rect 34928 66880 34936 66944
rect 35000 66896 35016 66944
rect 35080 66896 35096 66944
rect 35160 66896 35176 66944
rect 35240 66880 35248 66944
rect 34928 66660 34970 66880
rect 35206 66660 35248 66880
rect 34928 65856 35248 66660
rect 34928 65792 34936 65856
rect 35000 65792 35016 65856
rect 35080 65792 35096 65856
rect 35160 65792 35176 65856
rect 35240 65792 35248 65856
rect 34928 64768 35248 65792
rect 34928 64704 34936 64768
rect 35000 64704 35016 64768
rect 35080 64704 35096 64768
rect 35160 64704 35176 64768
rect 35240 64704 35248 64768
rect 34928 63680 35248 64704
rect 34928 63616 34936 63680
rect 35000 63616 35016 63680
rect 35080 63616 35096 63680
rect 35160 63616 35176 63680
rect 35240 63616 35248 63680
rect 34928 62592 35248 63616
rect 35588 101216 35908 101776
rect 35588 101152 35596 101216
rect 35660 101152 35676 101216
rect 35740 101152 35756 101216
rect 35820 101152 35836 101216
rect 35900 101152 35908 101216
rect 35588 100128 35908 101152
rect 35588 100064 35596 100128
rect 35660 100064 35676 100128
rect 35740 100064 35756 100128
rect 35820 100064 35836 100128
rect 35900 100064 35908 100128
rect 35588 99040 35908 100064
rect 35588 98976 35596 99040
rect 35660 98976 35676 99040
rect 35740 98976 35756 99040
rect 35820 98976 35836 99040
rect 35900 98976 35908 99040
rect 35588 98192 35908 98976
rect 35588 97956 35630 98192
rect 35866 97956 35908 98192
rect 35588 97952 35908 97956
rect 35588 97888 35596 97952
rect 35660 97888 35676 97952
rect 35740 97888 35756 97952
rect 35820 97888 35836 97952
rect 35900 97888 35908 97952
rect 35588 96864 35908 97888
rect 35588 96800 35596 96864
rect 35660 96800 35676 96864
rect 35740 96800 35756 96864
rect 35820 96800 35836 96864
rect 35900 96800 35908 96864
rect 35588 95776 35908 96800
rect 35588 95712 35596 95776
rect 35660 95712 35676 95776
rect 35740 95712 35756 95776
rect 35820 95712 35836 95776
rect 35900 95712 35908 95776
rect 35588 94688 35908 95712
rect 35588 94624 35596 94688
rect 35660 94624 35676 94688
rect 35740 94624 35756 94688
rect 35820 94624 35836 94688
rect 35900 94624 35908 94688
rect 35588 93600 35908 94624
rect 35588 93536 35596 93600
rect 35660 93536 35676 93600
rect 35740 93536 35756 93600
rect 35820 93536 35836 93600
rect 35900 93536 35908 93600
rect 35588 92512 35908 93536
rect 35588 92448 35596 92512
rect 35660 92448 35676 92512
rect 35740 92448 35756 92512
rect 35820 92448 35836 92512
rect 35900 92448 35908 92512
rect 35588 91424 35908 92448
rect 35588 91360 35596 91424
rect 35660 91360 35676 91424
rect 35740 91360 35756 91424
rect 35820 91360 35836 91424
rect 35900 91360 35908 91424
rect 35588 90336 35908 91360
rect 35588 90272 35596 90336
rect 35660 90272 35676 90336
rect 35740 90272 35756 90336
rect 35820 90272 35836 90336
rect 35900 90272 35908 90336
rect 35588 89248 35908 90272
rect 35588 89184 35596 89248
rect 35660 89184 35676 89248
rect 35740 89184 35756 89248
rect 35820 89184 35836 89248
rect 35900 89184 35908 89248
rect 35588 88160 35908 89184
rect 35588 88096 35596 88160
rect 35660 88096 35676 88160
rect 35740 88096 35756 88160
rect 35820 88096 35836 88160
rect 35900 88096 35908 88160
rect 35588 87072 35908 88096
rect 35588 87008 35596 87072
rect 35660 87008 35676 87072
rect 35740 87008 35756 87072
rect 35820 87008 35836 87072
rect 35900 87008 35908 87072
rect 35588 85984 35908 87008
rect 35588 85920 35596 85984
rect 35660 85920 35676 85984
rect 35740 85920 35756 85984
rect 35820 85920 35836 85984
rect 35900 85920 35908 85984
rect 35588 84896 35908 85920
rect 35588 84832 35596 84896
rect 35660 84832 35676 84896
rect 35740 84832 35756 84896
rect 35820 84832 35836 84896
rect 35900 84832 35908 84896
rect 35588 83808 35908 84832
rect 35588 83744 35596 83808
rect 35660 83744 35676 83808
rect 35740 83744 35756 83808
rect 35820 83744 35836 83808
rect 35900 83744 35908 83808
rect 35588 82720 35908 83744
rect 35588 82656 35596 82720
rect 35660 82656 35676 82720
rect 35740 82656 35756 82720
rect 35820 82656 35836 82720
rect 35900 82656 35908 82720
rect 35588 81632 35908 82656
rect 35588 81568 35596 81632
rect 35660 81568 35676 81632
rect 35740 81568 35756 81632
rect 35820 81568 35836 81632
rect 35900 81568 35908 81632
rect 35588 80544 35908 81568
rect 35588 80480 35596 80544
rect 35660 80480 35676 80544
rect 35740 80480 35756 80544
rect 35820 80480 35836 80544
rect 35900 80480 35908 80544
rect 35588 79456 35908 80480
rect 35588 79392 35596 79456
rect 35660 79392 35676 79456
rect 35740 79392 35756 79456
rect 35820 79392 35836 79456
rect 35900 79392 35908 79456
rect 35588 78368 35908 79392
rect 35588 78304 35596 78368
rect 35660 78304 35676 78368
rect 35740 78304 35756 78368
rect 35820 78304 35836 78368
rect 35900 78304 35908 78368
rect 35588 77280 35908 78304
rect 35588 77216 35596 77280
rect 35660 77216 35676 77280
rect 35740 77216 35756 77280
rect 35820 77216 35836 77280
rect 35900 77216 35908 77280
rect 35588 76192 35908 77216
rect 65648 101760 65968 101776
rect 65648 101696 65656 101760
rect 65720 101696 65736 101760
rect 65800 101696 65816 101760
rect 65880 101696 65896 101760
rect 65960 101696 65968 101760
rect 65648 100672 65968 101696
rect 65648 100608 65656 100672
rect 65720 100608 65736 100672
rect 65800 100608 65816 100672
rect 65880 100608 65896 100672
rect 65960 100608 65968 100672
rect 65648 99584 65968 100608
rect 65648 99520 65656 99584
rect 65720 99520 65736 99584
rect 65800 99520 65816 99584
rect 65880 99520 65896 99584
rect 65960 99520 65968 99584
rect 65648 98496 65968 99520
rect 65648 98432 65656 98496
rect 65720 98432 65736 98496
rect 65800 98432 65816 98496
rect 65880 98432 65896 98496
rect 65960 98432 65968 98496
rect 65648 97532 65968 98432
rect 65648 97408 65690 97532
rect 65926 97408 65968 97532
rect 65648 97344 65656 97408
rect 65960 97344 65968 97408
rect 65648 97296 65690 97344
rect 65926 97296 65968 97344
rect 65648 96320 65968 97296
rect 65648 96256 65656 96320
rect 65720 96256 65736 96320
rect 65800 96256 65816 96320
rect 65880 96256 65896 96320
rect 65960 96256 65968 96320
rect 65648 95232 65968 96256
rect 65648 95168 65656 95232
rect 65720 95168 65736 95232
rect 65800 95168 65816 95232
rect 65880 95168 65896 95232
rect 65960 95168 65968 95232
rect 65648 94144 65968 95168
rect 65648 94080 65656 94144
rect 65720 94080 65736 94144
rect 65800 94080 65816 94144
rect 65880 94080 65896 94144
rect 65960 94080 65968 94144
rect 65648 93056 65968 94080
rect 65648 92992 65656 93056
rect 65720 92992 65736 93056
rect 65800 92992 65816 93056
rect 65880 92992 65896 93056
rect 65960 92992 65968 93056
rect 65648 91968 65968 92992
rect 65648 91904 65656 91968
rect 65720 91904 65736 91968
rect 65800 91904 65816 91968
rect 65880 91904 65896 91968
rect 65960 91904 65968 91968
rect 65648 90880 65968 91904
rect 65648 90816 65656 90880
rect 65720 90816 65736 90880
rect 65800 90816 65816 90880
rect 65880 90816 65896 90880
rect 65960 90816 65968 90880
rect 65648 89792 65968 90816
rect 65648 89728 65656 89792
rect 65720 89728 65736 89792
rect 65800 89728 65816 89792
rect 65880 89728 65896 89792
rect 65960 89728 65968 89792
rect 65648 88704 65968 89728
rect 65648 88640 65656 88704
rect 65720 88640 65736 88704
rect 65800 88640 65816 88704
rect 65880 88640 65896 88704
rect 65960 88640 65968 88704
rect 65648 87616 65968 88640
rect 65648 87552 65656 87616
rect 65720 87552 65736 87616
rect 65800 87552 65816 87616
rect 65880 87552 65896 87616
rect 65960 87552 65968 87616
rect 65648 86528 65968 87552
rect 65648 86464 65656 86528
rect 65720 86464 65736 86528
rect 65800 86464 65816 86528
rect 65880 86464 65896 86528
rect 65960 86464 65968 86528
rect 65648 85440 65968 86464
rect 65648 85376 65656 85440
rect 65720 85376 65736 85440
rect 65800 85376 65816 85440
rect 65880 85376 65896 85440
rect 65960 85376 65968 85440
rect 65648 84352 65968 85376
rect 65648 84288 65656 84352
rect 65720 84288 65736 84352
rect 65800 84288 65816 84352
rect 65880 84288 65896 84352
rect 65960 84288 65968 84352
rect 65648 83264 65968 84288
rect 65648 83200 65656 83264
rect 65720 83200 65736 83264
rect 65800 83200 65816 83264
rect 65880 83200 65896 83264
rect 65960 83200 65968 83264
rect 65648 82176 65968 83200
rect 65648 82112 65656 82176
rect 65720 82112 65736 82176
rect 65800 82112 65816 82176
rect 65880 82112 65896 82176
rect 65960 82112 65968 82176
rect 65648 81088 65968 82112
rect 65648 81024 65656 81088
rect 65720 81024 65736 81088
rect 65800 81024 65816 81088
rect 65880 81024 65896 81088
rect 65960 81024 65968 81088
rect 65648 80000 65968 81024
rect 65648 79936 65656 80000
rect 65720 79936 65736 80000
rect 65800 79936 65816 80000
rect 65880 79936 65896 80000
rect 65960 79936 65968 80000
rect 65648 78912 65968 79936
rect 65648 78848 65656 78912
rect 65720 78848 65736 78912
rect 65800 78848 65816 78912
rect 65880 78848 65896 78912
rect 65960 78848 65968 78912
rect 65648 77824 65968 78848
rect 65648 77760 65656 77824
rect 65720 77760 65736 77824
rect 65800 77760 65816 77824
rect 65880 77760 65896 77824
rect 65960 77760 65968 77824
rect 45139 77076 45205 77077
rect 45139 77012 45140 77076
rect 45204 77012 45205 77076
rect 45139 77011 45205 77012
rect 37595 76260 37661 76261
rect 37595 76196 37596 76260
rect 37660 76196 37661 76260
rect 37595 76195 37661 76196
rect 35588 76128 35596 76192
rect 35660 76128 35676 76192
rect 35740 76128 35756 76192
rect 35820 76128 35836 76192
rect 35900 76128 35908 76192
rect 35588 75104 35908 76128
rect 35588 75040 35596 75104
rect 35660 75040 35676 75104
rect 35740 75040 35756 75104
rect 35820 75040 35836 75104
rect 35900 75040 35908 75104
rect 35588 74016 35908 75040
rect 35588 73952 35596 74016
rect 35660 73952 35676 74016
rect 35740 73952 35756 74016
rect 35820 73952 35836 74016
rect 35900 73952 35908 74016
rect 35588 72928 35908 73952
rect 35588 72864 35596 72928
rect 35660 72864 35676 72928
rect 35740 72864 35756 72928
rect 35820 72864 35836 72928
rect 35900 72864 35908 72928
rect 35588 71840 35908 72864
rect 35588 71776 35596 71840
rect 35660 71776 35676 71840
rect 35740 71776 35756 71840
rect 35820 71776 35836 71840
rect 35900 71776 35908 71840
rect 35588 70752 35908 71776
rect 35588 70688 35596 70752
rect 35660 70688 35676 70752
rect 35740 70688 35756 70752
rect 35820 70688 35836 70752
rect 35900 70688 35908 70752
rect 35588 69664 35908 70688
rect 35588 69600 35596 69664
rect 35660 69600 35676 69664
rect 35740 69600 35756 69664
rect 35820 69600 35836 69664
rect 35900 69600 35908 69664
rect 35588 68576 35908 69600
rect 35588 68512 35596 68576
rect 35660 68512 35676 68576
rect 35740 68512 35756 68576
rect 35820 68512 35836 68576
rect 35900 68512 35908 68576
rect 35588 67556 35908 68512
rect 35588 67488 35630 67556
rect 35866 67488 35908 67556
rect 35588 67424 35596 67488
rect 35900 67424 35908 67488
rect 35588 67320 35630 67424
rect 35866 67320 35908 67424
rect 35588 66400 35908 67320
rect 35588 66336 35596 66400
rect 35660 66336 35676 66400
rect 35740 66336 35756 66400
rect 35820 66336 35836 66400
rect 35900 66336 35908 66400
rect 35588 65312 35908 66336
rect 35588 65248 35596 65312
rect 35660 65248 35676 65312
rect 35740 65248 35756 65312
rect 35820 65248 35836 65312
rect 35900 65248 35908 65312
rect 35588 64224 35908 65248
rect 35588 64160 35596 64224
rect 35660 64160 35676 64224
rect 35740 64160 35756 64224
rect 35820 64160 35836 64224
rect 35900 64160 35908 64224
rect 35588 63136 35908 64160
rect 35588 63072 35596 63136
rect 35660 63072 35676 63136
rect 35740 63072 35756 63136
rect 35820 63072 35836 63136
rect 35900 63072 35908 63136
rect 35387 62796 35453 62797
rect 35387 62732 35388 62796
rect 35452 62732 35453 62796
rect 35387 62731 35453 62732
rect 34928 62528 34936 62592
rect 35000 62528 35016 62592
rect 35080 62528 35096 62592
rect 35160 62528 35176 62592
rect 35240 62528 35248 62592
rect 34928 61504 35248 62528
rect 34928 61440 34936 61504
rect 35000 61440 35016 61504
rect 35080 61440 35096 61504
rect 35160 61440 35176 61504
rect 35240 61440 35248 61504
rect 34928 60416 35248 61440
rect 34928 60352 34936 60416
rect 35000 60352 35016 60416
rect 35080 60352 35096 60416
rect 35160 60352 35176 60416
rect 35240 60352 35248 60416
rect 34928 59834 35248 60352
rect 4868 59650 5188 59808
rect 1668 58720 1676 58784
rect 1740 58720 1756 58784
rect 1820 58720 1828 58784
rect 1668 57696 1828 58720
rect 32570 58172 32636 58173
rect 32570 58108 32571 58172
rect 32635 58108 32636 58172
rect 35390 58170 35450 62731
rect 35588 62048 35908 63072
rect 35588 61984 35596 62048
rect 35660 61984 35676 62048
rect 35740 61984 35756 62048
rect 35820 61984 35836 62048
rect 35900 61984 35908 62048
rect 35588 60960 35908 61984
rect 35588 60896 35596 60960
rect 35660 60896 35676 60960
rect 35740 60896 35756 60960
rect 35820 60896 35836 60960
rect 35900 60896 35908 60960
rect 35588 59872 35908 60896
rect 35588 59808 35596 59872
rect 35660 59808 35676 59872
rect 35740 59808 35756 59872
rect 35820 59808 35836 59872
rect 35900 59808 35908 59872
rect 35588 59650 35908 59808
rect 37598 58170 37658 76195
rect 42563 75988 42629 75989
rect 42563 75924 42564 75988
rect 42628 75924 42629 75988
rect 42563 75923 42629 75924
rect 40171 74628 40237 74629
rect 40171 74564 40172 74628
rect 40236 74564 40237 74628
rect 40171 74563 40237 74564
rect 40174 58170 40234 74563
rect 32570 58107 32636 58108
rect 35069 58110 35450 58170
rect 37565 58110 37658 58170
rect 40082 58110 40234 58170
rect 30074 57900 30140 57901
rect 30074 57836 30075 57900
rect 30139 57836 30140 57900
rect 30074 57835 30140 57836
rect 1668 57632 1676 57696
rect 1740 57632 1756 57696
rect 1820 57632 1828 57696
rect 30077 57676 30137 57835
rect 32573 57676 32633 58107
rect 35069 57676 35129 58110
rect 37565 57676 37625 58110
rect 40082 57676 40142 58110
rect 42566 57676 42626 75923
rect 45142 58170 45202 77011
rect 65648 76736 65968 77760
rect 65648 76672 65656 76736
rect 65720 76672 65736 76736
rect 65800 76672 65816 76736
rect 65880 76672 65896 76736
rect 65960 76672 65968 76736
rect 50107 75852 50173 75853
rect 50107 75788 50108 75852
rect 50172 75788 50173 75852
rect 50107 75787 50173 75788
rect 47531 71908 47597 71909
rect 47531 71844 47532 71908
rect 47596 71844 47597 71908
rect 47531 71843 47597 71844
rect 45053 58110 45202 58170
rect 45053 57676 45113 58110
rect 47534 57676 47594 71843
rect 50110 58170 50170 75787
rect 65648 75648 65968 76672
rect 65648 75584 65656 75648
rect 65720 75584 65736 75648
rect 65800 75584 65816 75648
rect 65880 75584 65896 75648
rect 65960 75584 65968 75648
rect 52499 74628 52565 74629
rect 52499 74564 52500 74628
rect 52564 74564 52565 74628
rect 52499 74563 52565 74564
rect 50045 58110 50170 58170
rect 52502 58170 52562 74563
rect 65648 74560 65968 75584
rect 65648 74496 65656 74560
rect 65720 74496 65736 74560
rect 65800 74496 65816 74560
rect 65880 74496 65896 74560
rect 65960 74496 65968 74560
rect 55075 73948 55141 73949
rect 55075 73884 55076 73948
rect 55140 73884 55141 73948
rect 55075 73883 55141 73884
rect 55078 58170 55138 73883
rect 65648 73472 65968 74496
rect 65648 73408 65656 73472
rect 65720 73408 65736 73472
rect 65800 73408 65816 73472
rect 65880 73408 65896 73472
rect 65960 73408 65968 73472
rect 65648 72384 65968 73408
rect 65648 72320 65656 72384
rect 65720 72320 65736 72384
rect 65800 72320 65816 72384
rect 65880 72320 65896 72384
rect 65960 72320 65968 72384
rect 65648 71296 65968 72320
rect 65648 71232 65656 71296
rect 65720 71232 65736 71296
rect 65800 71232 65816 71296
rect 65880 71232 65896 71296
rect 65960 71232 65968 71296
rect 65648 70208 65968 71232
rect 65648 70144 65656 70208
rect 65720 70144 65736 70208
rect 65800 70144 65816 70208
rect 65880 70144 65896 70208
rect 65960 70144 65968 70208
rect 65648 69120 65968 70144
rect 65648 69056 65656 69120
rect 65720 69056 65736 69120
rect 65800 69056 65816 69120
rect 65880 69056 65896 69120
rect 65960 69056 65968 69120
rect 65648 68032 65968 69056
rect 65648 67968 65656 68032
rect 65720 67968 65736 68032
rect 65800 67968 65816 68032
rect 65880 67968 65896 68032
rect 65960 67968 65968 68032
rect 65648 66944 65968 67968
rect 65648 66880 65656 66944
rect 65720 66896 65736 66944
rect 65800 66896 65816 66944
rect 65880 66896 65896 66944
rect 65960 66880 65968 66944
rect 65648 66660 65690 66880
rect 65926 66660 65968 66880
rect 65648 65856 65968 66660
rect 65648 65792 65656 65856
rect 65720 65792 65736 65856
rect 65800 65792 65816 65856
rect 65880 65792 65896 65856
rect 65960 65792 65968 65856
rect 65648 64768 65968 65792
rect 65648 64704 65656 64768
rect 65720 64704 65736 64768
rect 65800 64704 65816 64768
rect 65880 64704 65896 64768
rect 65960 64704 65968 64768
rect 65648 63680 65968 64704
rect 65648 63616 65656 63680
rect 65720 63616 65736 63680
rect 65800 63616 65816 63680
rect 65880 63616 65896 63680
rect 65960 63616 65968 63680
rect 65648 62592 65968 63616
rect 65648 62528 65656 62592
rect 65720 62528 65736 62592
rect 65800 62528 65816 62592
rect 65880 62528 65896 62592
rect 65960 62528 65968 62592
rect 65648 61504 65968 62528
rect 65648 61440 65656 61504
rect 65720 61440 65736 61504
rect 65800 61440 65816 61504
rect 65880 61440 65896 61504
rect 65960 61440 65968 61504
rect 65648 60416 65968 61440
rect 65648 60352 65656 60416
rect 65720 60352 65736 60416
rect 65800 60352 65816 60416
rect 65880 60352 65896 60416
rect 65960 60352 65968 60416
rect 65648 59650 65968 60352
rect 66308 101216 66628 101776
rect 66308 101152 66316 101216
rect 66380 101152 66396 101216
rect 66460 101152 66476 101216
rect 66540 101152 66556 101216
rect 66620 101152 66628 101216
rect 66308 100128 66628 101152
rect 66308 100064 66316 100128
rect 66380 100064 66396 100128
rect 66460 100064 66476 100128
rect 66540 100064 66556 100128
rect 66620 100064 66628 100128
rect 66308 99040 66628 100064
rect 66308 98976 66316 99040
rect 66380 98976 66396 99040
rect 66460 98976 66476 99040
rect 66540 98976 66556 99040
rect 66620 98976 66628 99040
rect 66308 98192 66628 98976
rect 66308 97956 66350 98192
rect 66586 97956 66628 98192
rect 66308 97952 66628 97956
rect 66308 97888 66316 97952
rect 66380 97888 66396 97952
rect 66460 97888 66476 97952
rect 66540 97888 66556 97952
rect 66620 97888 66628 97952
rect 66308 96864 66628 97888
rect 66308 96800 66316 96864
rect 66380 96800 66396 96864
rect 66460 96800 66476 96864
rect 66540 96800 66556 96864
rect 66620 96800 66628 96864
rect 66308 95776 66628 96800
rect 66308 95712 66316 95776
rect 66380 95712 66396 95776
rect 66460 95712 66476 95776
rect 66540 95712 66556 95776
rect 66620 95712 66628 95776
rect 66308 94688 66628 95712
rect 66308 94624 66316 94688
rect 66380 94624 66396 94688
rect 66460 94624 66476 94688
rect 66540 94624 66556 94688
rect 66620 94624 66628 94688
rect 66308 93600 66628 94624
rect 66308 93536 66316 93600
rect 66380 93536 66396 93600
rect 66460 93536 66476 93600
rect 66540 93536 66556 93600
rect 66620 93536 66628 93600
rect 66308 92512 66628 93536
rect 66308 92448 66316 92512
rect 66380 92448 66396 92512
rect 66460 92448 66476 92512
rect 66540 92448 66556 92512
rect 66620 92448 66628 92512
rect 66308 91424 66628 92448
rect 66308 91360 66316 91424
rect 66380 91360 66396 91424
rect 66460 91360 66476 91424
rect 66540 91360 66556 91424
rect 66620 91360 66628 91424
rect 66308 90336 66628 91360
rect 66308 90272 66316 90336
rect 66380 90272 66396 90336
rect 66460 90272 66476 90336
rect 66540 90272 66556 90336
rect 66620 90272 66628 90336
rect 66308 89248 66628 90272
rect 66308 89184 66316 89248
rect 66380 89184 66396 89248
rect 66460 89184 66476 89248
rect 66540 89184 66556 89248
rect 66620 89184 66628 89248
rect 66308 88160 66628 89184
rect 66308 88096 66316 88160
rect 66380 88096 66396 88160
rect 66460 88096 66476 88160
rect 66540 88096 66556 88160
rect 66620 88096 66628 88160
rect 66308 87072 66628 88096
rect 66308 87008 66316 87072
rect 66380 87008 66396 87072
rect 66460 87008 66476 87072
rect 66540 87008 66556 87072
rect 66620 87008 66628 87072
rect 66308 85984 66628 87008
rect 66308 85920 66316 85984
rect 66380 85920 66396 85984
rect 66460 85920 66476 85984
rect 66540 85920 66556 85984
rect 66620 85920 66628 85984
rect 66308 84896 66628 85920
rect 66308 84832 66316 84896
rect 66380 84832 66396 84896
rect 66460 84832 66476 84896
rect 66540 84832 66556 84896
rect 66620 84832 66628 84896
rect 66308 83808 66628 84832
rect 66308 83744 66316 83808
rect 66380 83744 66396 83808
rect 66460 83744 66476 83808
rect 66540 83744 66556 83808
rect 66620 83744 66628 83808
rect 66308 82720 66628 83744
rect 66308 82656 66316 82720
rect 66380 82656 66396 82720
rect 66460 82656 66476 82720
rect 66540 82656 66556 82720
rect 66620 82656 66628 82720
rect 66308 81632 66628 82656
rect 66308 81568 66316 81632
rect 66380 81568 66396 81632
rect 66460 81568 66476 81632
rect 66540 81568 66556 81632
rect 66620 81568 66628 81632
rect 66308 80544 66628 81568
rect 66308 80480 66316 80544
rect 66380 80480 66396 80544
rect 66460 80480 66476 80544
rect 66540 80480 66556 80544
rect 66620 80480 66628 80544
rect 66308 79456 66628 80480
rect 66308 79392 66316 79456
rect 66380 79392 66396 79456
rect 66460 79392 66476 79456
rect 66540 79392 66556 79456
rect 66620 79392 66628 79456
rect 66308 78368 66628 79392
rect 66308 78304 66316 78368
rect 66380 78304 66396 78368
rect 66460 78304 66476 78368
rect 66540 78304 66556 78368
rect 66620 78304 66628 78368
rect 66308 77280 66628 78304
rect 66308 77216 66316 77280
rect 66380 77216 66396 77280
rect 66460 77216 66476 77280
rect 66540 77216 66556 77280
rect 66620 77216 66628 77280
rect 66308 76192 66628 77216
rect 66308 76128 66316 76192
rect 66380 76128 66396 76192
rect 66460 76128 66476 76192
rect 66540 76128 66556 76192
rect 66620 76128 66628 76192
rect 66308 75104 66628 76128
rect 66308 75040 66316 75104
rect 66380 75040 66396 75104
rect 66460 75040 66476 75104
rect 66540 75040 66556 75104
rect 66620 75040 66628 75104
rect 66308 74016 66628 75040
rect 66308 73952 66316 74016
rect 66380 73952 66396 74016
rect 66460 73952 66476 74016
rect 66540 73952 66556 74016
rect 66620 73952 66628 74016
rect 66308 72928 66628 73952
rect 66308 72864 66316 72928
rect 66380 72864 66396 72928
rect 66460 72864 66476 72928
rect 66540 72864 66556 72928
rect 66620 72864 66628 72928
rect 66308 71840 66628 72864
rect 66308 71776 66316 71840
rect 66380 71776 66396 71840
rect 66460 71776 66476 71840
rect 66540 71776 66556 71840
rect 66620 71776 66628 71840
rect 66308 70752 66628 71776
rect 66308 70688 66316 70752
rect 66380 70688 66396 70752
rect 66460 70688 66476 70752
rect 66540 70688 66556 70752
rect 66620 70688 66628 70752
rect 66308 69664 66628 70688
rect 66308 69600 66316 69664
rect 66380 69600 66396 69664
rect 66460 69600 66476 69664
rect 66540 69600 66556 69664
rect 66620 69600 66628 69664
rect 66308 68576 66628 69600
rect 66308 68512 66316 68576
rect 66380 68512 66396 68576
rect 66460 68512 66476 68576
rect 66540 68512 66556 68576
rect 66620 68512 66628 68576
rect 66308 67556 66628 68512
rect 66308 67488 66350 67556
rect 66586 67488 66628 67556
rect 66308 67424 66316 67488
rect 66620 67424 66628 67488
rect 66308 67320 66350 67424
rect 66586 67320 66628 67424
rect 66308 66400 66628 67320
rect 66308 66336 66316 66400
rect 66380 66336 66396 66400
rect 66460 66336 66476 66400
rect 66540 66336 66556 66400
rect 66620 66336 66628 66400
rect 66308 65312 66628 66336
rect 66308 65248 66316 65312
rect 66380 65248 66396 65312
rect 66460 65248 66476 65312
rect 66540 65248 66556 65312
rect 66620 65248 66628 65312
rect 66308 64224 66628 65248
rect 66308 64160 66316 64224
rect 66380 64160 66396 64224
rect 66460 64160 66476 64224
rect 66540 64160 66556 64224
rect 66620 64160 66628 64224
rect 66308 63136 66628 64160
rect 66308 63072 66316 63136
rect 66380 63072 66396 63136
rect 66460 63072 66476 63136
rect 66540 63072 66556 63136
rect 66620 63072 66628 63136
rect 66308 62048 66628 63072
rect 66308 61984 66316 62048
rect 66380 61984 66396 62048
rect 66460 61984 66476 62048
rect 66540 61984 66556 62048
rect 66620 61984 66628 62048
rect 66308 60960 66628 61984
rect 66308 60896 66316 60960
rect 66380 60896 66396 60960
rect 66460 60896 66476 60960
rect 66540 60896 66556 60960
rect 66620 60896 66628 60960
rect 66308 59872 66628 60896
rect 96368 101760 96688 101776
rect 96368 101696 96376 101760
rect 96440 101696 96456 101760
rect 96520 101696 96536 101760
rect 96600 101696 96616 101760
rect 96680 101696 96688 101760
rect 96368 100672 96688 101696
rect 96368 100608 96376 100672
rect 96440 100608 96456 100672
rect 96520 100608 96536 100672
rect 96600 100608 96616 100672
rect 96680 100608 96688 100672
rect 96368 99584 96688 100608
rect 96368 99520 96376 99584
rect 96440 99520 96456 99584
rect 96520 99520 96536 99584
rect 96600 99520 96616 99584
rect 96680 99520 96688 99584
rect 96368 98496 96688 99520
rect 96368 98432 96376 98496
rect 96440 98432 96456 98496
rect 96520 98432 96536 98496
rect 96600 98432 96616 98496
rect 96680 98432 96688 98496
rect 96368 97532 96688 98432
rect 96368 97408 96410 97532
rect 96646 97408 96688 97532
rect 96368 97344 96376 97408
rect 96680 97344 96688 97408
rect 96368 97296 96410 97344
rect 96646 97296 96688 97344
rect 96368 96320 96688 97296
rect 96368 96256 96376 96320
rect 96440 96256 96456 96320
rect 96520 96256 96536 96320
rect 96600 96256 96616 96320
rect 96680 96256 96688 96320
rect 96368 95232 96688 96256
rect 96368 95168 96376 95232
rect 96440 95168 96456 95232
rect 96520 95168 96536 95232
rect 96600 95168 96616 95232
rect 96680 95168 96688 95232
rect 96368 94144 96688 95168
rect 96368 94080 96376 94144
rect 96440 94080 96456 94144
rect 96520 94080 96536 94144
rect 96600 94080 96616 94144
rect 96680 94080 96688 94144
rect 96368 93056 96688 94080
rect 96368 92992 96376 93056
rect 96440 92992 96456 93056
rect 96520 92992 96536 93056
rect 96600 92992 96616 93056
rect 96680 92992 96688 93056
rect 96368 91968 96688 92992
rect 96368 91904 96376 91968
rect 96440 91904 96456 91968
rect 96520 91904 96536 91968
rect 96600 91904 96616 91968
rect 96680 91904 96688 91968
rect 96368 90880 96688 91904
rect 96368 90816 96376 90880
rect 96440 90816 96456 90880
rect 96520 90816 96536 90880
rect 96600 90816 96616 90880
rect 96680 90816 96688 90880
rect 96368 89792 96688 90816
rect 96368 89728 96376 89792
rect 96440 89728 96456 89792
rect 96520 89728 96536 89792
rect 96600 89728 96616 89792
rect 96680 89728 96688 89792
rect 96368 88704 96688 89728
rect 96368 88640 96376 88704
rect 96440 88640 96456 88704
rect 96520 88640 96536 88704
rect 96600 88640 96616 88704
rect 96680 88640 96688 88704
rect 96368 87616 96688 88640
rect 96368 87552 96376 87616
rect 96440 87552 96456 87616
rect 96520 87552 96536 87616
rect 96600 87552 96616 87616
rect 96680 87552 96688 87616
rect 96368 86528 96688 87552
rect 96368 86464 96376 86528
rect 96440 86464 96456 86528
rect 96520 86464 96536 86528
rect 96600 86464 96616 86528
rect 96680 86464 96688 86528
rect 96368 85440 96688 86464
rect 96368 85376 96376 85440
rect 96440 85376 96456 85440
rect 96520 85376 96536 85440
rect 96600 85376 96616 85440
rect 96680 85376 96688 85440
rect 96368 84352 96688 85376
rect 96368 84288 96376 84352
rect 96440 84288 96456 84352
rect 96520 84288 96536 84352
rect 96600 84288 96616 84352
rect 96680 84288 96688 84352
rect 96368 83264 96688 84288
rect 96368 83200 96376 83264
rect 96440 83200 96456 83264
rect 96520 83200 96536 83264
rect 96600 83200 96616 83264
rect 96680 83200 96688 83264
rect 96368 82176 96688 83200
rect 96368 82112 96376 82176
rect 96440 82112 96456 82176
rect 96520 82112 96536 82176
rect 96600 82112 96616 82176
rect 96680 82112 96688 82176
rect 96368 81088 96688 82112
rect 96368 81024 96376 81088
rect 96440 81024 96456 81088
rect 96520 81024 96536 81088
rect 96600 81024 96616 81088
rect 96680 81024 96688 81088
rect 96368 80000 96688 81024
rect 96368 79936 96376 80000
rect 96440 79936 96456 80000
rect 96520 79936 96536 80000
rect 96600 79936 96616 80000
rect 96680 79936 96688 80000
rect 96368 78912 96688 79936
rect 96368 78848 96376 78912
rect 96440 78848 96456 78912
rect 96520 78848 96536 78912
rect 96600 78848 96616 78912
rect 96680 78848 96688 78912
rect 96368 77824 96688 78848
rect 96368 77760 96376 77824
rect 96440 77760 96456 77824
rect 96520 77760 96536 77824
rect 96600 77760 96616 77824
rect 96680 77760 96688 77824
rect 96368 76736 96688 77760
rect 96368 76672 96376 76736
rect 96440 76672 96456 76736
rect 96520 76672 96536 76736
rect 96600 76672 96616 76736
rect 96680 76672 96688 76736
rect 96368 75648 96688 76672
rect 96368 75584 96376 75648
rect 96440 75584 96456 75648
rect 96520 75584 96536 75648
rect 96600 75584 96616 75648
rect 96680 75584 96688 75648
rect 96368 74560 96688 75584
rect 96368 74496 96376 74560
rect 96440 74496 96456 74560
rect 96520 74496 96536 74560
rect 96600 74496 96616 74560
rect 96680 74496 96688 74560
rect 96368 73472 96688 74496
rect 96368 73408 96376 73472
rect 96440 73408 96456 73472
rect 96520 73408 96536 73472
rect 96600 73408 96616 73472
rect 96680 73408 96688 73472
rect 96368 72384 96688 73408
rect 96368 72320 96376 72384
rect 96440 72320 96456 72384
rect 96520 72320 96536 72384
rect 96600 72320 96616 72384
rect 96680 72320 96688 72384
rect 96368 71296 96688 72320
rect 96368 71232 96376 71296
rect 96440 71232 96456 71296
rect 96520 71232 96536 71296
rect 96600 71232 96616 71296
rect 96680 71232 96688 71296
rect 96368 70208 96688 71232
rect 96368 70144 96376 70208
rect 96440 70144 96456 70208
rect 96520 70144 96536 70208
rect 96600 70144 96616 70208
rect 96680 70144 96688 70208
rect 96368 69120 96688 70144
rect 96368 69056 96376 69120
rect 96440 69056 96456 69120
rect 96520 69056 96536 69120
rect 96600 69056 96616 69120
rect 96680 69056 96688 69120
rect 96368 68032 96688 69056
rect 96368 67968 96376 68032
rect 96440 67968 96456 68032
rect 96520 67968 96536 68032
rect 96600 67968 96616 68032
rect 96680 67968 96688 68032
rect 96368 66944 96688 67968
rect 96368 66880 96376 66944
rect 96440 66896 96456 66944
rect 96520 66896 96536 66944
rect 96600 66896 96616 66944
rect 96680 66880 96688 66944
rect 96368 66660 96410 66880
rect 96646 66660 96688 66880
rect 96368 65856 96688 66660
rect 96368 65792 96376 65856
rect 96440 65792 96456 65856
rect 96520 65792 96536 65856
rect 96600 65792 96616 65856
rect 96680 65792 96688 65856
rect 96368 64768 96688 65792
rect 96368 64704 96376 64768
rect 96440 64704 96456 64768
rect 96520 64704 96536 64768
rect 96600 64704 96616 64768
rect 96680 64704 96688 64768
rect 96368 63680 96688 64704
rect 96368 63616 96376 63680
rect 96440 63616 96456 63680
rect 96520 63616 96536 63680
rect 96600 63616 96616 63680
rect 96680 63616 96688 63680
rect 96368 62592 96688 63616
rect 96368 62528 96376 62592
rect 96440 62528 96456 62592
rect 96520 62528 96536 62592
rect 96600 62528 96616 62592
rect 96680 62528 96688 62592
rect 96368 61504 96688 62528
rect 96368 61440 96376 61504
rect 96440 61440 96456 61504
rect 96520 61440 96536 61504
rect 96600 61440 96616 61504
rect 96680 61440 96688 61504
rect 67587 60756 67653 60757
rect 67587 60692 67588 60756
rect 67652 60692 67653 60756
rect 67587 60691 67653 60692
rect 66308 59808 66316 59872
rect 66380 59808 66396 59872
rect 66460 59808 66476 59872
rect 66540 59808 66556 59872
rect 66620 59808 66628 59872
rect 66308 59650 66628 59808
rect 57467 58852 57533 58853
rect 57467 58788 57468 58852
rect 57532 58788 57533 58852
rect 57467 58787 57533 58788
rect 52502 58110 52601 58170
rect 50045 57676 50105 58110
rect 52541 57676 52601 58110
rect 55037 58110 55138 58170
rect 57470 58170 57530 58787
rect 62619 58716 62685 58717
rect 62619 58652 62620 58716
rect 62684 58652 62685 58716
rect 62619 58651 62685 58652
rect 60043 58580 60109 58581
rect 60043 58516 60044 58580
rect 60108 58516 60109 58580
rect 60043 58515 60109 58516
rect 57470 58110 57593 58170
rect 55037 57676 55097 58110
rect 57533 57676 57593 58110
rect 60046 57676 60106 58515
rect 62622 58170 62682 58651
rect 67590 58170 67650 60691
rect 96368 60416 96688 61440
rect 96368 60352 96376 60416
rect 96440 60352 96456 60416
rect 96520 60352 96536 60416
rect 96600 60352 96616 60416
rect 96680 60352 96688 60416
rect 96368 59650 96688 60352
rect 97028 101216 97348 101776
rect 97028 101152 97036 101216
rect 97100 101152 97116 101216
rect 97180 101152 97196 101216
rect 97260 101152 97276 101216
rect 97340 101152 97348 101216
rect 97028 100128 97348 101152
rect 97028 100064 97036 100128
rect 97100 100064 97116 100128
rect 97180 100064 97196 100128
rect 97260 100064 97276 100128
rect 97340 100064 97348 100128
rect 97028 99040 97348 100064
rect 97028 98976 97036 99040
rect 97100 98976 97116 99040
rect 97180 98976 97196 99040
rect 97260 98976 97276 99040
rect 97340 98976 97348 99040
rect 97028 98192 97348 98976
rect 97028 97956 97070 98192
rect 97306 97956 97348 98192
rect 97028 97952 97348 97956
rect 97028 97888 97036 97952
rect 97100 97888 97116 97952
rect 97180 97888 97196 97952
rect 97260 97888 97276 97952
rect 97340 97888 97348 97952
rect 97028 96864 97348 97888
rect 97028 96800 97036 96864
rect 97100 96800 97116 96864
rect 97180 96800 97196 96864
rect 97260 96800 97276 96864
rect 97340 96800 97348 96864
rect 97028 95776 97348 96800
rect 97028 95712 97036 95776
rect 97100 95712 97116 95776
rect 97180 95712 97196 95776
rect 97260 95712 97276 95776
rect 97340 95712 97348 95776
rect 97028 94688 97348 95712
rect 97028 94624 97036 94688
rect 97100 94624 97116 94688
rect 97180 94624 97196 94688
rect 97260 94624 97276 94688
rect 97340 94624 97348 94688
rect 97028 93600 97348 94624
rect 97028 93536 97036 93600
rect 97100 93536 97116 93600
rect 97180 93536 97196 93600
rect 97260 93536 97276 93600
rect 97340 93536 97348 93600
rect 97028 92512 97348 93536
rect 97028 92448 97036 92512
rect 97100 92448 97116 92512
rect 97180 92448 97196 92512
rect 97260 92448 97276 92512
rect 97340 92448 97348 92512
rect 97028 91424 97348 92448
rect 97028 91360 97036 91424
rect 97100 91360 97116 91424
rect 97180 91360 97196 91424
rect 97260 91360 97276 91424
rect 97340 91360 97348 91424
rect 97028 90336 97348 91360
rect 97028 90272 97036 90336
rect 97100 90272 97116 90336
rect 97180 90272 97196 90336
rect 97260 90272 97276 90336
rect 97340 90272 97348 90336
rect 97028 89248 97348 90272
rect 97028 89184 97036 89248
rect 97100 89184 97116 89248
rect 97180 89184 97196 89248
rect 97260 89184 97276 89248
rect 97340 89184 97348 89248
rect 97028 88160 97348 89184
rect 97028 88096 97036 88160
rect 97100 88096 97116 88160
rect 97180 88096 97196 88160
rect 97260 88096 97276 88160
rect 97340 88096 97348 88160
rect 97028 87072 97348 88096
rect 97028 87008 97036 87072
rect 97100 87008 97116 87072
rect 97180 87008 97196 87072
rect 97260 87008 97276 87072
rect 97340 87008 97348 87072
rect 97028 85984 97348 87008
rect 97028 85920 97036 85984
rect 97100 85920 97116 85984
rect 97180 85920 97196 85984
rect 97260 85920 97276 85984
rect 97340 85920 97348 85984
rect 97028 84896 97348 85920
rect 97028 84832 97036 84896
rect 97100 84832 97116 84896
rect 97180 84832 97196 84896
rect 97260 84832 97276 84896
rect 97340 84832 97348 84896
rect 97028 83808 97348 84832
rect 97028 83744 97036 83808
rect 97100 83744 97116 83808
rect 97180 83744 97196 83808
rect 97260 83744 97276 83808
rect 97340 83744 97348 83808
rect 97028 82720 97348 83744
rect 97028 82656 97036 82720
rect 97100 82656 97116 82720
rect 97180 82656 97196 82720
rect 97260 82656 97276 82720
rect 97340 82656 97348 82720
rect 97028 81632 97348 82656
rect 97028 81568 97036 81632
rect 97100 81568 97116 81632
rect 97180 81568 97196 81632
rect 97260 81568 97276 81632
rect 97340 81568 97348 81632
rect 97028 80544 97348 81568
rect 97028 80480 97036 80544
rect 97100 80480 97116 80544
rect 97180 80480 97196 80544
rect 97260 80480 97276 80544
rect 97340 80480 97348 80544
rect 97028 79456 97348 80480
rect 97028 79392 97036 79456
rect 97100 79392 97116 79456
rect 97180 79392 97196 79456
rect 97260 79392 97276 79456
rect 97340 79392 97348 79456
rect 97028 78368 97348 79392
rect 97028 78304 97036 78368
rect 97100 78304 97116 78368
rect 97180 78304 97196 78368
rect 97260 78304 97276 78368
rect 97340 78304 97348 78368
rect 97028 77280 97348 78304
rect 97028 77216 97036 77280
rect 97100 77216 97116 77280
rect 97180 77216 97196 77280
rect 97260 77216 97276 77280
rect 97340 77216 97348 77280
rect 97028 76192 97348 77216
rect 97028 76128 97036 76192
rect 97100 76128 97116 76192
rect 97180 76128 97196 76192
rect 97260 76128 97276 76192
rect 97340 76128 97348 76192
rect 97028 75104 97348 76128
rect 97028 75040 97036 75104
rect 97100 75040 97116 75104
rect 97180 75040 97196 75104
rect 97260 75040 97276 75104
rect 97340 75040 97348 75104
rect 97028 74016 97348 75040
rect 97028 73952 97036 74016
rect 97100 73952 97116 74016
rect 97180 73952 97196 74016
rect 97260 73952 97276 74016
rect 97340 73952 97348 74016
rect 97028 72928 97348 73952
rect 97028 72864 97036 72928
rect 97100 72864 97116 72928
rect 97180 72864 97196 72928
rect 97260 72864 97276 72928
rect 97340 72864 97348 72928
rect 97028 71840 97348 72864
rect 97028 71776 97036 71840
rect 97100 71776 97116 71840
rect 97180 71776 97196 71840
rect 97260 71776 97276 71840
rect 97340 71776 97348 71840
rect 97028 70752 97348 71776
rect 97028 70688 97036 70752
rect 97100 70688 97116 70752
rect 97180 70688 97196 70752
rect 97260 70688 97276 70752
rect 97340 70688 97348 70752
rect 97028 69664 97348 70688
rect 97028 69600 97036 69664
rect 97100 69600 97116 69664
rect 97180 69600 97196 69664
rect 97260 69600 97276 69664
rect 97340 69600 97348 69664
rect 97028 68576 97348 69600
rect 97028 68512 97036 68576
rect 97100 68512 97116 68576
rect 97180 68512 97196 68576
rect 97260 68512 97276 68576
rect 97340 68512 97348 68576
rect 97028 67556 97348 68512
rect 97028 67488 97070 67556
rect 97306 67488 97348 67556
rect 97028 67424 97036 67488
rect 97340 67424 97348 67488
rect 97028 67320 97070 67424
rect 97306 67320 97348 67424
rect 97028 66400 97348 67320
rect 97028 66336 97036 66400
rect 97100 66336 97116 66400
rect 97180 66336 97196 66400
rect 97260 66336 97276 66400
rect 97340 66336 97348 66400
rect 97028 65312 97348 66336
rect 97028 65248 97036 65312
rect 97100 65248 97116 65312
rect 97180 65248 97196 65312
rect 97260 65248 97276 65312
rect 97340 65248 97348 65312
rect 97028 64224 97348 65248
rect 97028 64160 97036 64224
rect 97100 64160 97116 64224
rect 97180 64160 97196 64224
rect 97260 64160 97276 64224
rect 97340 64160 97348 64224
rect 97028 63136 97348 64160
rect 97028 63072 97036 63136
rect 97100 63072 97116 63136
rect 97180 63072 97196 63136
rect 97260 63072 97276 63136
rect 97340 63072 97348 63136
rect 97028 62048 97348 63072
rect 97028 61984 97036 62048
rect 97100 61984 97116 62048
rect 97180 61984 97196 62048
rect 97260 61984 97276 62048
rect 97340 61984 97348 62048
rect 97028 60960 97348 61984
rect 97028 60896 97036 60960
rect 97100 60896 97116 60960
rect 97180 60896 97196 60960
rect 97260 60896 97276 60960
rect 97340 60896 97348 60960
rect 97028 59872 97348 60896
rect 97028 59808 97036 59872
rect 97100 59808 97116 59872
rect 97180 59808 97196 59872
rect 97260 59808 97276 59872
rect 97340 59808 97348 59872
rect 97028 59650 97348 59808
rect 98924 60416 99244 60432
rect 98924 60352 98932 60416
rect 98996 60352 99012 60416
rect 99076 60352 99092 60416
rect 99156 60352 99172 60416
rect 99236 60352 99244 60416
rect 98924 59328 99244 60352
rect 98924 59264 98932 59328
rect 98996 59264 99012 59328
rect 99076 59264 99092 59328
rect 99156 59264 99172 59328
rect 99236 59264 99244 59328
rect 98924 58240 99244 59264
rect 98924 58176 98932 58240
rect 98996 58176 99012 58240
rect 99076 58176 99092 58240
rect 99156 58176 99172 58240
rect 99236 58176 99244 58240
rect 62530 58110 62682 58170
rect 67517 58110 67650 58170
rect 80141 58172 80207 58173
rect 62530 57676 62590 58110
rect 65018 57900 65084 57901
rect 65018 57836 65019 57900
rect 65083 57836 65084 57900
rect 65018 57835 65084 57836
rect 65021 57676 65081 57835
rect 67517 57676 67577 58110
rect 80141 58108 80142 58172
rect 80206 58108 80207 58172
rect 80141 58107 80207 58108
rect 80144 57676 80204 58107
rect 81309 58036 81375 58037
rect 81309 57972 81310 58036
rect 81374 57972 81375 58036
rect 81309 57971 81375 57972
rect 81312 57676 81372 57971
rect 89857 57900 89923 57901
rect 89857 57836 89858 57900
rect 89922 57836 89923 57900
rect 89857 57835 89923 57836
rect 89860 57676 89920 57835
rect 1668 56608 1828 57632
rect 1668 56544 1676 56608
rect 1740 56544 1756 56608
rect 1820 56544 1828 56608
rect 1668 55520 1828 56544
rect 1668 55456 1676 55520
rect 1740 55456 1756 55520
rect 1820 55456 1828 55520
rect 1668 54432 1828 55456
rect 1668 54368 1676 54432
rect 1740 54368 1756 54432
rect 1820 54368 1828 54432
rect 1668 53344 1828 54368
rect 1668 53280 1676 53344
rect 1740 53280 1756 53344
rect 1820 53280 1828 53344
rect 1668 52256 1828 53280
rect 1668 52192 1676 52256
rect 1740 52192 1756 52256
rect 1820 52192 1828 52256
rect 1668 51168 1828 52192
rect 1668 51104 1676 51168
rect 1740 51104 1756 51168
rect 1820 51104 1828 51168
rect 1668 50080 1828 51104
rect 1668 50016 1676 50080
rect 1740 50016 1756 50080
rect 1820 50016 1828 50080
rect 1668 48992 1828 50016
rect 1668 48928 1676 48992
rect 1740 48928 1756 48992
rect 1820 48928 1828 48992
rect 1668 47904 1828 48928
rect 1668 47840 1676 47904
rect 1740 47840 1756 47904
rect 1820 47840 1828 47904
rect 1668 46816 1828 47840
rect 1668 46752 1676 46816
rect 1740 46752 1756 46816
rect 1820 46752 1828 46816
rect 1668 45728 1828 46752
rect 1668 45664 1676 45728
rect 1740 45664 1756 45728
rect 1820 45664 1828 45728
rect 1668 44640 1828 45664
rect 1668 44576 1676 44640
rect 1740 44576 1756 44640
rect 1820 44576 1828 44640
rect 1668 43552 1828 44576
rect 1668 43488 1676 43552
rect 1740 43488 1756 43552
rect 1820 43488 1828 43552
rect 1668 42464 1828 43488
rect 1668 42400 1676 42464
rect 1740 42400 1756 42464
rect 1820 42400 1828 42464
rect 1668 41376 1828 42400
rect 1668 41312 1676 41376
rect 1740 41312 1756 41376
rect 1820 41312 1828 41376
rect 1668 40288 1828 41312
rect 1668 40224 1676 40288
rect 1740 40224 1756 40288
rect 1820 40224 1828 40288
rect 1668 39200 1828 40224
rect 1668 39136 1676 39200
rect 1740 39136 1756 39200
rect 1820 39136 1828 39200
rect 1668 38112 1828 39136
rect 1668 38048 1676 38112
rect 1740 38048 1756 38112
rect 1820 38048 1828 38112
rect 1668 37024 1828 38048
rect 1668 36960 1676 37024
rect 1740 36960 1756 37024
rect 1820 36960 1828 37024
rect 98924 57152 99244 58176
rect 98924 57088 98932 57152
rect 98996 57088 99012 57152
rect 99076 57088 99092 57152
rect 99156 57088 99172 57152
rect 99236 57088 99244 57152
rect 98924 56064 99244 57088
rect 98924 56000 98932 56064
rect 98996 56000 99012 56064
rect 99076 56000 99092 56064
rect 99156 56000 99172 56064
rect 99236 56000 99244 56064
rect 98924 54976 99244 56000
rect 98924 54912 98932 54976
rect 98996 54912 99012 54976
rect 99076 54912 99092 54976
rect 99156 54912 99172 54976
rect 99236 54912 99244 54976
rect 98924 53888 99244 54912
rect 98924 53824 98932 53888
rect 98996 53824 99012 53888
rect 99076 53824 99092 53888
rect 99156 53824 99172 53888
rect 99236 53824 99244 53888
rect 98924 52800 99244 53824
rect 98924 52736 98932 52800
rect 98996 52736 99012 52800
rect 99076 52736 99092 52800
rect 99156 52736 99172 52800
rect 99236 52736 99244 52800
rect 98924 51712 99244 52736
rect 98924 51648 98932 51712
rect 98996 51648 99012 51712
rect 99076 51648 99092 51712
rect 99156 51648 99172 51712
rect 99236 51648 99244 51712
rect 98924 50624 99244 51648
rect 98924 50560 98932 50624
rect 98996 50560 99012 50624
rect 99076 50560 99092 50624
rect 99156 50560 99172 50624
rect 99236 50560 99244 50624
rect 98924 49536 99244 50560
rect 98924 49472 98932 49536
rect 98996 49472 99012 49536
rect 99076 49472 99092 49536
rect 99156 49472 99172 49536
rect 99236 49472 99244 49536
rect 98924 48448 99244 49472
rect 98924 48384 98932 48448
rect 98996 48384 99012 48448
rect 99076 48384 99092 48448
rect 99156 48384 99172 48448
rect 99236 48384 99244 48448
rect 98924 47360 99244 48384
rect 98924 47296 98932 47360
rect 98996 47296 99012 47360
rect 99076 47296 99092 47360
rect 99156 47296 99172 47360
rect 99236 47296 99244 47360
rect 98924 46272 99244 47296
rect 98924 46208 98932 46272
rect 98996 46208 99012 46272
rect 99076 46208 99092 46272
rect 99156 46208 99172 46272
rect 99236 46208 99244 46272
rect 98924 45184 99244 46208
rect 98924 45120 98932 45184
rect 98996 45120 99012 45184
rect 99076 45120 99092 45184
rect 99156 45120 99172 45184
rect 99236 45120 99244 45184
rect 98924 44096 99244 45120
rect 98924 44032 98932 44096
rect 98996 44032 99012 44096
rect 99076 44032 99092 44096
rect 99156 44032 99172 44096
rect 99236 44032 99244 44096
rect 98924 43008 99244 44032
rect 98924 42944 98932 43008
rect 98996 42944 99012 43008
rect 99076 42944 99092 43008
rect 99156 42944 99172 43008
rect 99236 42944 99244 43008
rect 98924 41920 99244 42944
rect 98924 41856 98932 41920
rect 98996 41856 99012 41920
rect 99076 41856 99092 41920
rect 99156 41856 99172 41920
rect 99236 41856 99244 41920
rect 98924 40832 99244 41856
rect 98924 40768 98932 40832
rect 98996 40768 99012 40832
rect 99076 40768 99092 40832
rect 99156 40768 99172 40832
rect 99236 40768 99244 40832
rect 98924 39744 99244 40768
rect 98924 39680 98932 39744
rect 98996 39680 99012 39744
rect 99076 39680 99092 39744
rect 99156 39680 99172 39744
rect 99236 39680 99244 39744
rect 98924 38656 99244 39680
rect 98924 38592 98932 38656
rect 98996 38592 99012 38656
rect 99076 38592 99092 38656
rect 99156 38592 99172 38656
rect 99236 38592 99244 38656
rect 98924 37568 99244 38592
rect 98924 37504 98932 37568
rect 98996 37504 99012 37568
rect 99076 37504 99092 37568
rect 99156 37504 99172 37568
rect 99236 37504 99244 37568
rect 1668 35936 1828 36960
rect 4696 36920 5044 36962
rect 4696 36684 4752 36920
rect 4988 36684 5044 36920
rect 4696 36642 5044 36684
rect 94936 36920 95284 36962
rect 94936 36684 94992 36920
rect 95228 36684 95284 36920
rect 94936 36642 95284 36684
rect 98924 36480 99244 37504
rect 98924 36416 98932 36480
rect 98996 36416 99012 36480
rect 99076 36416 99092 36480
rect 99156 36416 99172 36480
rect 99236 36416 99244 36480
rect 4000 36260 4348 36302
rect 4000 36024 4056 36260
rect 4292 36024 4348 36260
rect 4000 35982 4348 36024
rect 95632 36260 95980 36302
rect 95632 36024 95688 36260
rect 95924 36024 95980 36260
rect 95632 35982 95980 36024
rect 98924 36260 99244 36416
rect 98924 36024 98966 36260
rect 99202 36024 99244 36260
rect 1668 35872 1676 35936
rect 1740 35872 1756 35936
rect 1820 35872 1828 35936
rect 1668 34848 1828 35872
rect 1668 34784 1676 34848
rect 1740 34784 1756 34848
rect 1820 34784 1828 34848
rect 1668 33760 1828 34784
rect 1668 33696 1676 33760
rect 1740 33696 1756 33760
rect 1820 33696 1828 33760
rect 1668 32672 1828 33696
rect 1668 32608 1676 32672
rect 1740 32608 1756 32672
rect 1820 32608 1828 32672
rect 1668 31584 1828 32608
rect 1668 31520 1676 31584
rect 1740 31520 1756 31584
rect 1820 31520 1828 31584
rect 1668 30496 1828 31520
rect 1668 30432 1676 30496
rect 1740 30432 1756 30496
rect 1820 30432 1828 30496
rect 1668 29408 1828 30432
rect 1668 29344 1676 29408
rect 1740 29344 1756 29408
rect 1820 29344 1828 29408
rect 1668 28320 1828 29344
rect 1668 28256 1676 28320
rect 1740 28256 1756 28320
rect 1820 28256 1828 28320
rect 1668 27232 1828 28256
rect 1668 27168 1676 27232
rect 1740 27168 1756 27232
rect 1820 27168 1828 27232
rect 1668 26144 1828 27168
rect 1668 26080 1676 26144
rect 1740 26080 1756 26144
rect 1820 26080 1828 26144
rect 1668 25056 1828 26080
rect 1668 24992 1676 25056
rect 1740 24992 1756 25056
rect 1820 24992 1828 25056
rect 1668 23968 1828 24992
rect 1668 23904 1676 23968
rect 1740 23904 1756 23968
rect 1820 23904 1828 23968
rect 1668 22880 1828 23904
rect 1668 22816 1676 22880
rect 1740 22816 1756 22880
rect 1820 22816 1828 22880
rect 1668 21792 1828 22816
rect 1668 21728 1676 21792
rect 1740 21728 1756 21792
rect 1820 21728 1828 21792
rect 1668 20704 1828 21728
rect 1668 20640 1676 20704
rect 1740 20640 1756 20704
rect 1820 20640 1828 20704
rect 1668 19616 1828 20640
rect 1668 19552 1676 19616
rect 1740 19552 1756 19616
rect 1820 19552 1828 19616
rect 1668 18528 1828 19552
rect 1668 18464 1676 18528
rect 1740 18464 1756 18528
rect 1820 18464 1828 18528
rect 1668 17440 1828 18464
rect 1668 17376 1676 17440
rect 1740 17376 1756 17440
rect 1820 17376 1828 17440
rect 1668 16352 1828 17376
rect 1668 16288 1676 16352
rect 1740 16288 1756 16352
rect 1820 16288 1828 16352
rect 1668 15264 1828 16288
rect 1668 15200 1676 15264
rect 1740 15200 1756 15264
rect 1820 15200 1828 15264
rect 1668 14176 1828 15200
rect 1668 14112 1676 14176
rect 1740 14112 1756 14176
rect 1820 14112 1828 14176
rect 1668 13088 1828 14112
rect 1668 13024 1676 13088
rect 1740 13024 1756 13088
rect 1820 13024 1828 13088
rect 1668 12000 1828 13024
rect 1668 11936 1676 12000
rect 1740 11936 1756 12000
rect 1820 11936 1828 12000
rect 1668 10912 1828 11936
rect 1668 10848 1676 10912
rect 1740 10848 1756 10912
rect 1820 10848 1828 10912
rect 1668 9824 1828 10848
rect 1668 9760 1676 9824
rect 1740 9760 1756 9824
rect 1820 9760 1828 9824
rect 1668 8736 1828 9760
rect 1668 8672 1676 8736
rect 1740 8672 1756 8736
rect 1820 8672 1828 8736
rect 1668 7648 1828 8672
rect 1668 7584 1676 7648
rect 1740 7584 1756 7648
rect 1820 7584 1828 7648
rect 1668 6560 1828 7584
rect 1668 6496 1676 6560
rect 1740 6496 1756 6560
rect 1820 6496 1828 6560
rect 1668 5472 1828 6496
rect 98924 35392 99244 36024
rect 98924 35328 98932 35392
rect 98996 35328 99012 35392
rect 99076 35328 99092 35392
rect 99156 35328 99172 35392
rect 99236 35328 99244 35392
rect 98924 34304 99244 35328
rect 98924 34240 98932 34304
rect 98996 34240 99012 34304
rect 99076 34240 99092 34304
rect 99156 34240 99172 34304
rect 99236 34240 99244 34304
rect 98924 33216 99244 34240
rect 98924 33152 98932 33216
rect 98996 33152 99012 33216
rect 99076 33152 99092 33216
rect 99156 33152 99172 33216
rect 99236 33152 99244 33216
rect 98924 32128 99244 33152
rect 98924 32064 98932 32128
rect 98996 32064 99012 32128
rect 99076 32064 99092 32128
rect 99156 32064 99172 32128
rect 99236 32064 99244 32128
rect 98924 31040 99244 32064
rect 98924 30976 98932 31040
rect 98996 30976 99012 31040
rect 99076 30976 99092 31040
rect 99156 30976 99172 31040
rect 99236 30976 99244 31040
rect 98924 29952 99244 30976
rect 98924 29888 98932 29952
rect 98996 29888 99012 29952
rect 99076 29888 99092 29952
rect 99156 29888 99172 29952
rect 99236 29888 99244 29952
rect 98924 28864 99244 29888
rect 98924 28800 98932 28864
rect 98996 28800 99012 28864
rect 99076 28800 99092 28864
rect 99156 28800 99172 28864
rect 99236 28800 99244 28864
rect 98924 27776 99244 28800
rect 98924 27712 98932 27776
rect 98996 27712 99012 27776
rect 99076 27712 99092 27776
rect 99156 27712 99172 27776
rect 99236 27712 99244 27776
rect 98924 26688 99244 27712
rect 98924 26624 98932 26688
rect 98996 26624 99012 26688
rect 99076 26624 99092 26688
rect 99156 26624 99172 26688
rect 99236 26624 99244 26688
rect 98924 25600 99244 26624
rect 98924 25536 98932 25600
rect 98996 25536 99012 25600
rect 99076 25536 99092 25600
rect 99156 25536 99172 25600
rect 99236 25536 99244 25600
rect 98924 24512 99244 25536
rect 98924 24448 98932 24512
rect 98996 24448 99012 24512
rect 99076 24448 99092 24512
rect 99156 24448 99172 24512
rect 99236 24448 99244 24512
rect 98924 23424 99244 24448
rect 98924 23360 98932 23424
rect 98996 23360 99012 23424
rect 99076 23360 99092 23424
rect 99156 23360 99172 23424
rect 99236 23360 99244 23424
rect 98924 22336 99244 23360
rect 98924 22272 98932 22336
rect 98996 22272 99012 22336
rect 99076 22272 99092 22336
rect 99156 22272 99172 22336
rect 99236 22272 99244 22336
rect 98924 21248 99244 22272
rect 98924 21184 98932 21248
rect 98996 21184 99012 21248
rect 99076 21184 99092 21248
rect 99156 21184 99172 21248
rect 99236 21184 99244 21248
rect 98924 20160 99244 21184
rect 98924 20096 98932 20160
rect 98996 20096 99012 20160
rect 99076 20096 99092 20160
rect 99156 20096 99172 20160
rect 99236 20096 99244 20160
rect 98924 19072 99244 20096
rect 98924 19008 98932 19072
rect 98996 19008 99012 19072
rect 99076 19008 99092 19072
rect 99156 19008 99172 19072
rect 99236 19008 99244 19072
rect 98924 17984 99244 19008
rect 98924 17920 98932 17984
rect 98996 17920 99012 17984
rect 99076 17920 99092 17984
rect 99156 17920 99172 17984
rect 99236 17920 99244 17984
rect 98924 16896 99244 17920
rect 98924 16832 98932 16896
rect 98996 16832 99012 16896
rect 99076 16832 99092 16896
rect 99156 16832 99172 16896
rect 99236 16832 99244 16896
rect 98924 15808 99244 16832
rect 98924 15744 98932 15808
rect 98996 15744 99012 15808
rect 99076 15744 99092 15808
rect 99156 15744 99172 15808
rect 99236 15744 99244 15808
rect 98924 14720 99244 15744
rect 98924 14656 98932 14720
rect 98996 14656 99012 14720
rect 99076 14656 99092 14720
rect 99156 14656 99172 14720
rect 99236 14656 99244 14720
rect 98924 13632 99244 14656
rect 98924 13568 98932 13632
rect 98996 13568 99012 13632
rect 99076 13568 99092 13632
rect 99156 13568 99172 13632
rect 99236 13568 99244 13632
rect 98924 12544 99244 13568
rect 98924 12480 98932 12544
rect 98996 12480 99012 12544
rect 99076 12480 99092 12544
rect 99156 12480 99172 12544
rect 99236 12480 99244 12544
rect 98924 11456 99244 12480
rect 98924 11392 98932 11456
rect 98996 11392 99012 11456
rect 99076 11392 99092 11456
rect 99156 11392 99172 11456
rect 99236 11392 99244 11456
rect 98924 10368 99244 11392
rect 98924 10304 98932 10368
rect 98996 10304 99012 10368
rect 99076 10304 99092 10368
rect 99156 10304 99172 10368
rect 99236 10304 99244 10368
rect 98924 9280 99244 10304
rect 98924 9216 98932 9280
rect 98996 9216 99012 9280
rect 99076 9216 99092 9280
rect 99156 9216 99172 9280
rect 99236 9216 99244 9280
rect 98924 8192 99244 9216
rect 98924 8128 98932 8192
rect 98996 8128 99012 8192
rect 99076 8128 99092 8192
rect 99156 8128 99172 8192
rect 99236 8128 99244 8192
rect 98924 7104 99244 8128
rect 98924 7040 98932 7104
rect 98996 7040 99012 7104
rect 99076 7040 99092 7104
rect 99156 7040 99172 7104
rect 99236 7040 99244 7104
rect 4696 6284 5044 6326
rect 4696 6048 4752 6284
rect 4988 6048 5044 6284
rect 4696 6006 5044 6048
rect 94936 6284 95284 6326
rect 94936 6048 94992 6284
rect 95228 6048 95284 6284
rect 94936 6006 95284 6048
rect 98924 6016 99244 7040
rect 98924 5952 98932 6016
rect 98996 5952 99012 6016
rect 99076 5952 99092 6016
rect 99156 5952 99172 6016
rect 99236 5952 99244 6016
rect 1668 5408 1676 5472
rect 1740 5408 1756 5472
rect 1820 5408 1828 5472
rect 1668 4384 1828 5408
rect 4000 5624 4348 5666
rect 4000 5388 4056 5624
rect 4292 5388 4348 5624
rect 4000 5346 4348 5388
rect 95632 5624 95980 5666
rect 95632 5388 95688 5624
rect 95924 5388 95980 5624
rect 95632 5346 95980 5388
rect 98924 5624 99244 5952
rect 98924 5388 98966 5624
rect 99202 5388 99244 5624
rect 1668 4320 1676 4384
rect 1740 4320 1756 4384
rect 1820 4320 1828 4384
rect 1668 3296 1828 4320
rect 98924 4928 99244 5388
rect 98924 4864 98932 4928
rect 98996 4864 99012 4928
rect 99076 4864 99092 4928
rect 99156 4864 99172 4928
rect 99236 4864 99244 4928
rect 10060 3909 10120 4038
rect 10057 3908 10123 3909
rect 10057 3844 10058 3908
rect 10122 3844 10123 3908
rect 10057 3843 10123 3844
rect 17440 3501 17500 4038
rect 18608 3770 18668 4038
rect 18608 3710 18706 3770
rect 17437 3500 17503 3501
rect 17437 3436 17438 3500
rect 17502 3436 17503 3500
rect 17437 3435 17503 3436
rect 1668 3232 1676 3296
rect 1740 3232 1756 3296
rect 1820 3232 1828 3296
rect 1668 2208 1828 3232
rect 18646 2821 18706 3710
rect 19776 3501 19836 4038
rect 20944 3501 21004 4038
rect 22112 3501 22172 4038
rect 23280 3770 23340 4038
rect 23246 3710 23340 3770
rect 19773 3500 19839 3501
rect 19773 3436 19774 3500
rect 19838 3436 19839 3500
rect 19773 3435 19839 3436
rect 20941 3500 21007 3501
rect 20941 3436 20942 3500
rect 21006 3436 21007 3500
rect 20941 3435 21007 3436
rect 22109 3500 22175 3501
rect 22109 3436 22110 3500
rect 22174 3436 22175 3500
rect 22109 3435 22175 3436
rect 23246 2821 23306 3710
rect 24448 3501 24508 4038
rect 25616 3501 25676 4038
rect 26784 3501 26844 4038
rect 27938 3501 27998 4038
rect 24445 3500 24511 3501
rect 24445 3436 24446 3500
rect 24510 3436 24511 3500
rect 24445 3435 24511 3436
rect 25613 3500 25679 3501
rect 25613 3436 25614 3500
rect 25678 3436 25679 3500
rect 25613 3435 25679 3436
rect 26781 3500 26847 3501
rect 26781 3436 26782 3500
rect 26846 3436 26847 3500
rect 26781 3435 26847 3436
rect 27935 3500 28001 3501
rect 27935 3436 27936 3500
rect 28000 3436 28001 3500
rect 27935 3435 28001 3436
rect 29134 2821 29194 4038
rect 30288 3501 30348 4038
rect 31456 3770 31516 4038
rect 31456 3710 31586 3770
rect 30285 3500 30351 3501
rect 30285 3436 30286 3500
rect 30350 3436 30351 3500
rect 30285 3435 30351 3436
rect 31526 2821 31586 3710
rect 32630 2821 32690 4038
rect 33792 3501 33852 4038
rect 34960 3501 35020 4038
rect 33789 3500 33855 3501
rect 33789 3436 33790 3500
rect 33854 3436 33855 3500
rect 33789 3435 33855 3436
rect 34957 3500 35023 3501
rect 34957 3436 34958 3500
rect 35022 3436 35023 3500
rect 34957 3435 35023 3436
rect 36126 2821 36186 4038
rect 37296 3770 37356 4038
rect 37230 3710 37356 3770
rect 37230 2821 37290 3710
rect 84529 3637 84589 4038
rect 84667 3773 84727 4038
rect 84816 3909 84876 4038
rect 84813 3908 84879 3909
rect 84813 3844 84814 3908
rect 84878 3844 84879 3908
rect 84813 3843 84879 3844
rect 98924 3840 99244 4864
rect 98924 3776 98932 3840
rect 98996 3776 99012 3840
rect 99076 3776 99092 3840
rect 99156 3776 99172 3840
rect 99236 3776 99244 3840
rect 84664 3772 84730 3773
rect 84664 3708 84665 3772
rect 84729 3708 84730 3772
rect 84664 3707 84730 3708
rect 84526 3636 84592 3637
rect 84526 3572 84527 3636
rect 84591 3572 84592 3636
rect 84526 3571 84592 3572
rect 18643 2820 18709 2821
rect 18643 2756 18644 2820
rect 18708 2756 18709 2820
rect 18643 2755 18709 2756
rect 23243 2820 23309 2821
rect 23243 2756 23244 2820
rect 23308 2756 23309 2820
rect 23243 2755 23309 2756
rect 29131 2820 29197 2821
rect 29131 2756 29132 2820
rect 29196 2756 29197 2820
rect 29131 2755 29197 2756
rect 31523 2820 31589 2821
rect 31523 2756 31524 2820
rect 31588 2756 31589 2820
rect 31523 2755 31589 2756
rect 32627 2820 32693 2821
rect 32627 2756 32628 2820
rect 32692 2756 32693 2820
rect 32627 2755 32693 2756
rect 36123 2820 36189 2821
rect 36123 2756 36124 2820
rect 36188 2756 36189 2820
rect 36123 2755 36189 2756
rect 37227 2820 37293 2821
rect 37227 2756 37228 2820
rect 37292 2756 37293 2820
rect 37227 2755 37293 2756
rect 1668 2144 1676 2208
rect 1740 2144 1756 2208
rect 1820 2144 1828 2208
rect 1668 2128 1828 2144
rect 98924 2752 99244 3776
rect 98924 2688 98932 2752
rect 98996 2688 99012 2752
rect 99076 2688 99092 2752
rect 99156 2688 99172 2752
rect 99236 2688 99244 2752
rect 98924 2128 99244 2688
rect 99660 59872 99980 60432
rect 99660 59808 99668 59872
rect 99732 59808 99748 59872
rect 99812 59808 99828 59872
rect 99892 59808 99908 59872
rect 99972 59808 99980 59872
rect 99660 58784 99980 59808
rect 99660 58720 99668 58784
rect 99732 58720 99748 58784
rect 99812 58720 99828 58784
rect 99892 58720 99908 58784
rect 99972 58720 99980 58784
rect 99660 57696 99980 58720
rect 99660 57632 99668 57696
rect 99732 57632 99748 57696
rect 99812 57632 99828 57696
rect 99892 57632 99908 57696
rect 99972 57632 99980 57696
rect 99660 56608 99980 57632
rect 99660 56544 99668 56608
rect 99732 56544 99748 56608
rect 99812 56544 99828 56608
rect 99892 56544 99908 56608
rect 99972 56544 99980 56608
rect 99660 55520 99980 56544
rect 99660 55456 99668 55520
rect 99732 55456 99748 55520
rect 99812 55456 99828 55520
rect 99892 55456 99908 55520
rect 99972 55456 99980 55520
rect 99660 54432 99980 55456
rect 99660 54368 99668 54432
rect 99732 54368 99748 54432
rect 99812 54368 99828 54432
rect 99892 54368 99908 54432
rect 99972 54368 99980 54432
rect 99660 53344 99980 54368
rect 99660 53280 99668 53344
rect 99732 53280 99748 53344
rect 99812 53280 99828 53344
rect 99892 53280 99908 53344
rect 99972 53280 99980 53344
rect 99660 52256 99980 53280
rect 99660 52192 99668 52256
rect 99732 52192 99748 52256
rect 99812 52192 99828 52256
rect 99892 52192 99908 52256
rect 99972 52192 99980 52256
rect 99660 51168 99980 52192
rect 99660 51104 99668 51168
rect 99732 51104 99748 51168
rect 99812 51104 99828 51168
rect 99892 51104 99908 51168
rect 99972 51104 99980 51168
rect 99660 50080 99980 51104
rect 99660 50016 99668 50080
rect 99732 50016 99748 50080
rect 99812 50016 99828 50080
rect 99892 50016 99908 50080
rect 99972 50016 99980 50080
rect 99660 48992 99980 50016
rect 99660 48928 99668 48992
rect 99732 48928 99748 48992
rect 99812 48928 99828 48992
rect 99892 48928 99908 48992
rect 99972 48928 99980 48992
rect 99660 47904 99980 48928
rect 99660 47840 99668 47904
rect 99732 47840 99748 47904
rect 99812 47840 99828 47904
rect 99892 47840 99908 47904
rect 99972 47840 99980 47904
rect 99660 46816 99980 47840
rect 99660 46752 99668 46816
rect 99732 46752 99748 46816
rect 99812 46752 99828 46816
rect 99892 46752 99908 46816
rect 99972 46752 99980 46816
rect 99660 45728 99980 46752
rect 99660 45664 99668 45728
rect 99732 45664 99748 45728
rect 99812 45664 99828 45728
rect 99892 45664 99908 45728
rect 99972 45664 99980 45728
rect 99660 44640 99980 45664
rect 99660 44576 99668 44640
rect 99732 44576 99748 44640
rect 99812 44576 99828 44640
rect 99892 44576 99908 44640
rect 99972 44576 99980 44640
rect 99660 43552 99980 44576
rect 99660 43488 99668 43552
rect 99732 43488 99748 43552
rect 99812 43488 99828 43552
rect 99892 43488 99908 43552
rect 99972 43488 99980 43552
rect 99660 42464 99980 43488
rect 99660 42400 99668 42464
rect 99732 42400 99748 42464
rect 99812 42400 99828 42464
rect 99892 42400 99908 42464
rect 99972 42400 99980 42464
rect 99660 41376 99980 42400
rect 99660 41312 99668 41376
rect 99732 41312 99748 41376
rect 99812 41312 99828 41376
rect 99892 41312 99908 41376
rect 99972 41312 99980 41376
rect 99660 40288 99980 41312
rect 99660 40224 99668 40288
rect 99732 40224 99748 40288
rect 99812 40224 99828 40288
rect 99892 40224 99908 40288
rect 99972 40224 99980 40288
rect 99660 39200 99980 40224
rect 99660 39136 99668 39200
rect 99732 39136 99748 39200
rect 99812 39136 99828 39200
rect 99892 39136 99908 39200
rect 99972 39136 99980 39200
rect 99660 38112 99980 39136
rect 99660 38048 99668 38112
rect 99732 38048 99748 38112
rect 99812 38048 99828 38112
rect 99892 38048 99908 38112
rect 99972 38048 99980 38112
rect 99660 37024 99980 38048
rect 99660 36960 99668 37024
rect 99732 36960 99748 37024
rect 99812 36960 99828 37024
rect 99892 36960 99908 37024
rect 99972 36960 99980 37024
rect 99660 36920 99980 36960
rect 99660 36684 99702 36920
rect 99938 36684 99980 36920
rect 99660 35936 99980 36684
rect 99660 35872 99668 35936
rect 99732 35872 99748 35936
rect 99812 35872 99828 35936
rect 99892 35872 99908 35936
rect 99972 35872 99980 35936
rect 99660 34848 99980 35872
rect 99660 34784 99668 34848
rect 99732 34784 99748 34848
rect 99812 34784 99828 34848
rect 99892 34784 99908 34848
rect 99972 34784 99980 34848
rect 99660 33760 99980 34784
rect 99660 33696 99668 33760
rect 99732 33696 99748 33760
rect 99812 33696 99828 33760
rect 99892 33696 99908 33760
rect 99972 33696 99980 33760
rect 99660 32672 99980 33696
rect 99660 32608 99668 32672
rect 99732 32608 99748 32672
rect 99812 32608 99828 32672
rect 99892 32608 99908 32672
rect 99972 32608 99980 32672
rect 99660 31584 99980 32608
rect 99660 31520 99668 31584
rect 99732 31520 99748 31584
rect 99812 31520 99828 31584
rect 99892 31520 99908 31584
rect 99972 31520 99980 31584
rect 99660 30496 99980 31520
rect 99660 30432 99668 30496
rect 99732 30432 99748 30496
rect 99812 30432 99828 30496
rect 99892 30432 99908 30496
rect 99972 30432 99980 30496
rect 99660 29408 99980 30432
rect 99660 29344 99668 29408
rect 99732 29344 99748 29408
rect 99812 29344 99828 29408
rect 99892 29344 99908 29408
rect 99972 29344 99980 29408
rect 99660 28320 99980 29344
rect 99660 28256 99668 28320
rect 99732 28256 99748 28320
rect 99812 28256 99828 28320
rect 99892 28256 99908 28320
rect 99972 28256 99980 28320
rect 99660 27232 99980 28256
rect 99660 27168 99668 27232
rect 99732 27168 99748 27232
rect 99812 27168 99828 27232
rect 99892 27168 99908 27232
rect 99972 27168 99980 27232
rect 99660 26144 99980 27168
rect 99660 26080 99668 26144
rect 99732 26080 99748 26144
rect 99812 26080 99828 26144
rect 99892 26080 99908 26144
rect 99972 26080 99980 26144
rect 99660 25056 99980 26080
rect 99660 24992 99668 25056
rect 99732 24992 99748 25056
rect 99812 24992 99828 25056
rect 99892 24992 99908 25056
rect 99972 24992 99980 25056
rect 99660 23968 99980 24992
rect 99660 23904 99668 23968
rect 99732 23904 99748 23968
rect 99812 23904 99828 23968
rect 99892 23904 99908 23968
rect 99972 23904 99980 23968
rect 99660 22880 99980 23904
rect 99660 22816 99668 22880
rect 99732 22816 99748 22880
rect 99812 22816 99828 22880
rect 99892 22816 99908 22880
rect 99972 22816 99980 22880
rect 99660 21792 99980 22816
rect 99660 21728 99668 21792
rect 99732 21728 99748 21792
rect 99812 21728 99828 21792
rect 99892 21728 99908 21792
rect 99972 21728 99980 21792
rect 99660 20704 99980 21728
rect 99660 20640 99668 20704
rect 99732 20640 99748 20704
rect 99812 20640 99828 20704
rect 99892 20640 99908 20704
rect 99972 20640 99980 20704
rect 99660 19616 99980 20640
rect 99660 19552 99668 19616
rect 99732 19552 99748 19616
rect 99812 19552 99828 19616
rect 99892 19552 99908 19616
rect 99972 19552 99980 19616
rect 99660 18528 99980 19552
rect 99660 18464 99668 18528
rect 99732 18464 99748 18528
rect 99812 18464 99828 18528
rect 99892 18464 99908 18528
rect 99972 18464 99980 18528
rect 99660 17440 99980 18464
rect 99660 17376 99668 17440
rect 99732 17376 99748 17440
rect 99812 17376 99828 17440
rect 99892 17376 99908 17440
rect 99972 17376 99980 17440
rect 99660 16352 99980 17376
rect 99660 16288 99668 16352
rect 99732 16288 99748 16352
rect 99812 16288 99828 16352
rect 99892 16288 99908 16352
rect 99972 16288 99980 16352
rect 99660 15264 99980 16288
rect 99660 15200 99668 15264
rect 99732 15200 99748 15264
rect 99812 15200 99828 15264
rect 99892 15200 99908 15264
rect 99972 15200 99980 15264
rect 99660 14176 99980 15200
rect 99660 14112 99668 14176
rect 99732 14112 99748 14176
rect 99812 14112 99828 14176
rect 99892 14112 99908 14176
rect 99972 14112 99980 14176
rect 99660 13088 99980 14112
rect 99660 13024 99668 13088
rect 99732 13024 99748 13088
rect 99812 13024 99828 13088
rect 99892 13024 99908 13088
rect 99972 13024 99980 13088
rect 99660 12000 99980 13024
rect 99660 11936 99668 12000
rect 99732 11936 99748 12000
rect 99812 11936 99828 12000
rect 99892 11936 99908 12000
rect 99972 11936 99980 12000
rect 99660 10912 99980 11936
rect 99660 10848 99668 10912
rect 99732 10848 99748 10912
rect 99812 10848 99828 10912
rect 99892 10848 99908 10912
rect 99972 10848 99980 10912
rect 99660 9824 99980 10848
rect 99660 9760 99668 9824
rect 99732 9760 99748 9824
rect 99812 9760 99828 9824
rect 99892 9760 99908 9824
rect 99972 9760 99980 9824
rect 99660 8736 99980 9760
rect 99660 8672 99668 8736
rect 99732 8672 99748 8736
rect 99812 8672 99828 8736
rect 99892 8672 99908 8736
rect 99972 8672 99980 8736
rect 99660 7648 99980 8672
rect 99660 7584 99668 7648
rect 99732 7584 99748 7648
rect 99812 7584 99828 7648
rect 99892 7584 99908 7648
rect 99972 7584 99980 7648
rect 99660 6560 99980 7584
rect 99660 6496 99668 6560
rect 99732 6496 99748 6560
rect 99812 6496 99828 6560
rect 99892 6496 99908 6560
rect 99972 6496 99980 6560
rect 99660 6284 99980 6496
rect 99660 6048 99702 6284
rect 99938 6048 99980 6284
rect 99660 5472 99980 6048
rect 99660 5408 99668 5472
rect 99732 5408 99748 5472
rect 99812 5408 99828 5472
rect 99892 5408 99908 5472
rect 99972 5408 99980 5472
rect 99660 4384 99980 5408
rect 99660 4320 99668 4384
rect 99732 4320 99748 4384
rect 99812 4320 99828 4384
rect 99892 4320 99908 4384
rect 99972 4320 99980 4384
rect 99660 3296 99980 4320
rect 99660 3232 99668 3296
rect 99732 3232 99748 3296
rect 99812 3232 99828 3296
rect 99892 3232 99908 3296
rect 99972 3232 99980 3296
rect 99660 2208 99980 3232
rect 99660 2144 99668 2208
rect 99732 2144 99748 2208
rect 99812 2144 99828 2208
rect 99892 2144 99908 2208
rect 99972 2144 99980 2208
rect 99660 2128 99980 2144
<< via4 >>
rect 4250 97408 4486 97532
rect 4250 97344 4280 97408
rect 4280 97344 4296 97408
rect 4296 97344 4360 97408
rect 4360 97344 4376 97408
rect 4376 97344 4440 97408
rect 4440 97344 4456 97408
rect 4456 97344 4486 97408
rect 4250 97296 4486 97344
rect 4250 66880 4280 66896
rect 4280 66880 4296 66896
rect 4296 66880 4360 66896
rect 4360 66880 4376 66896
rect 4376 66880 4440 66896
rect 4440 66880 4456 66896
rect 4456 66880 4486 66896
rect 4250 66660 4486 66880
rect 4910 97956 5146 98192
rect 4910 67488 5146 67556
rect 4910 67424 4940 67488
rect 4940 67424 4956 67488
rect 4956 67424 5020 67488
rect 5020 67424 5036 67488
rect 5036 67424 5100 67488
rect 5100 67424 5116 67488
rect 5116 67424 5146 67488
rect 4910 67320 5146 67424
rect 34970 97408 35206 97532
rect 34970 97344 35000 97408
rect 35000 97344 35016 97408
rect 35016 97344 35080 97408
rect 35080 97344 35096 97408
rect 35096 97344 35160 97408
rect 35160 97344 35176 97408
rect 35176 97344 35206 97408
rect 34970 97296 35206 97344
rect 34970 66880 35000 66896
rect 35000 66880 35016 66896
rect 35016 66880 35080 66896
rect 35080 66880 35096 66896
rect 35096 66880 35160 66896
rect 35160 66880 35176 66896
rect 35176 66880 35206 66896
rect 34970 66660 35206 66880
rect 35630 97956 35866 98192
rect 65690 97408 65926 97532
rect 65690 97344 65720 97408
rect 65720 97344 65736 97408
rect 65736 97344 65800 97408
rect 65800 97344 65816 97408
rect 65816 97344 65880 97408
rect 65880 97344 65896 97408
rect 65896 97344 65926 97408
rect 65690 97296 65926 97344
rect 35630 67488 35866 67556
rect 35630 67424 35660 67488
rect 35660 67424 35676 67488
rect 35676 67424 35740 67488
rect 35740 67424 35756 67488
rect 35756 67424 35820 67488
rect 35820 67424 35836 67488
rect 35836 67424 35866 67488
rect 35630 67320 35866 67424
rect 65690 66880 65720 66896
rect 65720 66880 65736 66896
rect 65736 66880 65800 66896
rect 65800 66880 65816 66896
rect 65816 66880 65880 66896
rect 65880 66880 65896 66896
rect 65896 66880 65926 66896
rect 65690 66660 65926 66880
rect 66350 97956 66586 98192
rect 66350 67488 66586 67556
rect 66350 67424 66380 67488
rect 66380 67424 66396 67488
rect 66396 67424 66460 67488
rect 66460 67424 66476 67488
rect 66476 67424 66540 67488
rect 66540 67424 66556 67488
rect 66556 67424 66586 67488
rect 66350 67320 66586 67424
rect 96410 97408 96646 97532
rect 96410 97344 96440 97408
rect 96440 97344 96456 97408
rect 96456 97344 96520 97408
rect 96520 97344 96536 97408
rect 96536 97344 96600 97408
rect 96600 97344 96616 97408
rect 96616 97344 96646 97408
rect 96410 97296 96646 97344
rect 96410 66880 96440 66896
rect 96440 66880 96456 66896
rect 96456 66880 96520 66896
rect 96520 66880 96536 66896
rect 96536 66880 96600 66896
rect 96600 66880 96616 66896
rect 96616 66880 96646 66896
rect 96410 66660 96646 66880
rect 97070 97956 97306 98192
rect 97070 67488 97306 67556
rect 97070 67424 97100 67488
rect 97100 67424 97116 67488
rect 97116 67424 97180 67488
rect 97180 67424 97196 67488
rect 97196 67424 97260 67488
rect 97260 67424 97276 67488
rect 97276 67424 97306 67488
rect 97070 67320 97306 67424
rect 4752 36684 4988 36920
rect 94992 36684 95228 36920
rect 4056 36024 4292 36260
rect 95688 36024 95924 36260
rect 98966 36024 99202 36260
rect 4752 6048 4988 6284
rect 94992 6048 95228 6284
rect 4056 5388 4292 5624
rect 95688 5388 95924 5624
rect 98966 5388 99202 5624
rect 99702 36684 99938 36920
rect 99702 6048 99938 6284
<< metal5 >>
rect 1056 98192 100880 98234
rect 1056 97956 4910 98192
rect 5146 97956 35630 98192
rect 35866 97956 66350 98192
rect 66586 97956 97070 98192
rect 97306 97956 100880 98192
rect 1056 97914 100880 97956
rect 1056 97532 100880 97574
rect 1056 97296 4250 97532
rect 4486 97296 34970 97532
rect 35206 97296 65690 97532
rect 65926 97296 96410 97532
rect 96646 97296 100880 97532
rect 1056 97254 100880 97296
rect 1056 67556 100880 67598
rect 1056 67320 4910 67556
rect 5146 67320 35630 67556
rect 35866 67320 66350 67556
rect 66586 67320 97070 67556
rect 97306 67320 100880 67556
rect 1056 67278 100880 67320
rect 1056 66896 100880 66938
rect 1056 66660 4250 66896
rect 4486 66660 34970 66896
rect 35206 66660 65690 66896
rect 65926 66660 96410 66896
rect 96646 66660 100880 66896
rect 1056 66618 100880 66660
rect 1056 36920 100880 36962
rect 1056 36684 4752 36920
rect 4988 36684 94992 36920
rect 95228 36684 99702 36920
rect 99938 36684 100880 36920
rect 1056 36642 100880 36684
rect 1056 36260 100880 36302
rect 1056 36024 4056 36260
rect 4292 36024 95688 36260
rect 95924 36024 98966 36260
rect 99202 36024 100880 36260
rect 1056 35982 100880 36024
rect 1056 6284 100880 6326
rect 1056 6048 4752 6284
rect 4988 6048 94992 6284
rect 95228 6048 99702 6284
rect 99938 6048 100880 6284
rect 1056 6006 100880 6048
rect 1056 5624 100880 5666
rect 1056 5388 4056 5624
rect 4292 5388 95688 5624
rect 95924 5388 98966 5624
rect 99202 5388 100880 5624
rect 1056 5346 100880 5388
use sky130_fd_sc_hd__inv_2  _040_
timestamp 1
transform 1 0 85836 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _041_
timestamp 1
transform -1 0 53360 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _042_
timestamp 1
transform -1 0 88320 0 1 59840
box -38 -48 682 592
use sky130_fd_sc_hd__and3_2  _043_
timestamp 1
transform 1 0 98256 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _044_
timestamp 1
transform -1 0 98624 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _045_
timestamp 1
transform -1 0 98532 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _046_
timestamp 1
transform -1 0 100004 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _047_
timestamp 1
transform -1 0 100188 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _048_
timestamp 1
transform -1 0 99820 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _049_
timestamp 1
transform 1 0 99084 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _050_
timestamp 1
transform 1 0 98256 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _051_
timestamp 1
transform -1 0 98992 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _052_
timestamp 1
transform 1 0 98256 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _053_
timestamp 1
transform -1 0 99084 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _054_
timestamp 1
transform -1 0 99544 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _055_
timestamp 1
transform 1 0 98256 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _056_
timestamp 1
transform -1 0 55016 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _057_
timestamp 1
transform -1 0 57040 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _058_
timestamp 1
transform -1 0 58512 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _059_
timestamp 1
transform 1 0 60536 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _060_
timestamp 1
transform -1 0 77280 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _061_
timestamp 1
transform 1 0 78476 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _062_
timestamp 1
transform 1 0 79212 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _063_
timestamp 1
transform 1 0 80132 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _064_
timestamp 1
transform 1 0 81696 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _065_
timestamp 1
transform 1 0 83904 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _066_
timestamp 1
transform 1 0 84364 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _067_
timestamp 1
transform 1 0 98256 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _068_
timestamp 1
transform 1 0 98256 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _069_
timestamp 1
transform 1 0 98256 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _070_
timestamp 1
transform 1 0 98256 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _071_
timestamp 1
transform 1 0 98348 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _072_
timestamp 1
transform 1 0 98348 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _073_
timestamp 1
transform -1 0 29348 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _074_
timestamp 1
transform -1 0 30544 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _075_
timestamp 1
transform -1 0 46736 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _076_
timestamp 1
transform -1 0 48392 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _077_
timestamp 1
transform -1 0 50140 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _078_
timestamp 1
transform -1 0 52072 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _079_
timestamp 1
transform 1 0 49404 0 -1 77248
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _080_
timestamp 1
transform 1 0 51336 0 1 77248
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _081_
timestamp 1
transform 1 0 53360 0 1 77248
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _082_
timestamp 1
transform 1 0 55568 0 1 77248
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _083_
timestamp 1
transform 1 0 57408 0 1 77248
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _084_
timestamp 1
transform 1 0 77004 0 1 60928
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _085_
timestamp 1
transform 1 0 78844 0 1 60928
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _086_
timestamp 1
transform 1 0 79672 0 -1 60928
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _087_
timestamp 1
transform 1 0 81512 0 -1 60928
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _088_
timestamp 1
transform 1 0 82064 0 1 60928
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _089_
timestamp 1
transform -1 0 86020 0 -1 60928
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _090_
timestamp 1
transform -1 0 87952 0 -1 60928
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _091_
timestamp 1
transform -1 0 100188 0 -1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _092_
timestamp 1
transform -1 0 100188 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _093_
timestamp 1
transform -1 0 100096 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _094_
timestamp 1
transform -1 0 100188 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _095_
timestamp 1
transform -1 0 100280 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _096_
timestamp 1
transform -1 0 100188 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _097_
timestamp 1
transform -1 0 22908 0 1 60928
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _098_
timestamp 1
transform -1 0 24380 0 -1 60928
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _099_
timestamp 1
transform 1 0 41768 0 1 77248
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _100_
timestamp 1
transform 1 0 43608 0 -1 77248
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _101_
timestamp 1
transform 1 0 45724 0 1 77248
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _102_
timestamp 1
transform 1 0 47932 0 1 77248
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1
transform 1 0 57408 0 -1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1
transform 1 0 76820 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1
transform -1 0 80868 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1
transform -1 0 79672 0 -1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1
transform -1 0 83536 0 -1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1
transform 1 0 81880 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1
transform 1 0 41768 0 -1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1
transform 1 0 41584 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1
transform 1 0 43608 0 1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1
transform 1 0 45724 0 -1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1
transform 1 0 47932 0 -1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1
transform 1 0 49404 0 1 76160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1
transform 1 0 51336 0 -1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1
transform 1 0 53360 0 -1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1
transform 1 0 55568 0 -1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1
transform -1 0 1932 0 1 62016
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1
transform 1 0 22356 0 -1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 1
transform -1 0 57132 0 1 59840
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1
transform -1 0 49956 0 1 59840
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1
transform 1 0 73692 0 1 59840
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkload0
timestamp 1
transform 1 0 48116 0 -1 60928
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_4  fanout18
timestamp 1
transform -1 0 60536 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  fanout19
timestamp 1
transform 1 0 98348 0 -1 26112
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_4  fanout20
timestamp 1
transform -1 0 98992 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3
timestamp 1
transform 1 0 1380 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1056
timestamp 1636968456
transform 1 0 98256 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1068
timestamp 1636968456
transform 1 0 99360 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1080
timestamp 1
transform 1 0 100464 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_3
timestamp 1
transform 1 0 1380 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1056
timestamp 1636968456
transform 1 0 98256 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_1068
timestamp 1636968456
transform 1 0 99360 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_1080
timestamp 1
transform 1 0 100464 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_3
timestamp 1
transform 1 0 1380 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1056
timestamp 1636968456
transform 1 0 98256 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_1068
timestamp 1636968456
transform 1 0 99360 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_1080
timestamp 1
transform 1 0 100464 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_3
timestamp 1
transform 1 0 1380 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1056
timestamp 1636968456
transform 1 0 98256 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_1068
timestamp 1636968456
transform 1 0 99360 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_1080
timestamp 1
transform 1 0 100464 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_3
timestamp 1
transform 1 0 1380 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1056
timestamp 1636968456
transform 1 0 98256 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_1068
timestamp 1636968456
transform 1 0 99360 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_1080
timestamp 1
transform 1 0 100464 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_3
timestamp 1
transform 1 0 1380 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1056
timestamp 1636968456
transform 1 0 98256 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_1068
timestamp 1636968456
transform 1 0 99360 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_1080
timestamp 1
transform 1 0 100464 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_3
timestamp 1
transform 1 0 1380 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1056
timestamp 1636968456
transform 1 0 98256 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_1068
timestamp 1636968456
transform 1 0 99360 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_1080
timestamp 1
transform 1 0 100464 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_3
timestamp 1
transform 1 0 1380 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1056
timestamp 1636968456
transform 1 0 98256 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_1068
timestamp 1636968456
transform 1 0 99360 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_1080
timestamp 1
transform 1 0 100464 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_3
timestamp 1
transform 1 0 1380 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1056
timestamp 1636968456
transform 1 0 98256 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_1068
timestamp 1636968456
transform 1 0 99360 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_1080
timestamp 1
transform 1 0 100464 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3
timestamp 1
transform 1 0 1380 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1056
timestamp 1636968456
transform 1 0 98256 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_1068
timestamp 1636968456
transform 1 0 99360 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_1080
timestamp 1
transform 1 0 100464 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_3
timestamp 1
transform 1 0 1380 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1056
timestamp 1636968456
transform 1 0 98256 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_1068
timestamp 1636968456
transform 1 0 99360 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_1080
timestamp 1
transform 1 0 100464 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_3
timestamp 1
transform 1 0 1380 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1056
timestamp 1636968456
transform 1 0 98256 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_1068
timestamp 1636968456
transform 1 0 99360 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_1080
timestamp 1
transform 1 0 100464 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_3
timestamp 1
transform 1 0 1380 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1056
timestamp 1636968456
transform 1 0 98256 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_1068
timestamp 1636968456
transform 1 0 99360 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_1080
timestamp 1
transform 1 0 100464 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_3
timestamp 1
transform 1 0 1380 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1056
timestamp 1636968456
transform 1 0 98256 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_1068
timestamp 1636968456
transform 1 0 99360 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_1080
timestamp 1
transform 1 0 100464 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_3
timestamp 1
transform 1 0 1380 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1056
timestamp 1636968456
transform 1 0 98256 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_1068
timestamp 1636968456
transform 1 0 99360 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_1080
timestamp 1
transform 1 0 100464 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_3
timestamp 1
transform 1 0 1380 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1056
timestamp 1636968456
transform 1 0 98256 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_1068
timestamp 1636968456
transform 1 0 99360 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_1080
timestamp 1
transform 1 0 100464 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_3
timestamp 1
transform 1 0 1380 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1056
timestamp 1636968456
transform 1 0 98256 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_1068
timestamp 1636968456
transform 1 0 99360 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_1080
timestamp 1
transform 1 0 100464 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_3
timestamp 1
transform 1 0 1380 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1056
timestamp 1636968456
transform 1 0 98256 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_1068
timestamp 1636968456
transform 1 0 99360 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_1080
timestamp 1
transform 1 0 100464 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_3
timestamp 1
transform 1 0 1380 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1056
timestamp 1636968456
transform 1 0 98256 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_1068
timestamp 1636968456
transform 1 0 99360 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_1080
timestamp 1
transform 1 0 100464 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_3
timestamp 1
transform 1 0 1380 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1056
timestamp 1636968456
transform 1 0 98256 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_1068
timestamp 1636968456
transform 1 0 99360 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_1080
timestamp 1
transform 1 0 100464 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_3
timestamp 1
transform 1 0 1380 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1056
timestamp 1636968456
transform 1 0 98256 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_1068
timestamp 1636968456
transform 1 0 99360 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_1080
timestamp 1
transform 1 0 100464 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_3
timestamp 1
transform 1 0 1380 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1056
timestamp 1636968456
transform 1 0 98256 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_1068
timestamp 1636968456
transform 1 0 99360 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_1080
timestamp 1
transform 1 0 100464 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_3
timestamp 1
transform 1 0 1380 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1056
timestamp 1636968456
transform 1 0 98256 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_1068
timestamp 1636968456
transform 1 0 99360 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_1080
timestamp 1
transform 1 0 100464 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_3
timestamp 1
transform 1 0 1380 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1056
timestamp 1636968456
transform 1 0 98256 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_1068
timestamp 1636968456
transform 1 0 99360 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_1080
timestamp 1
transform 1 0 100464 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_3
timestamp 1
transform 1 0 1380 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1056
timestamp 1636968456
transform 1 0 98256 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_1068
timestamp 1636968456
transform 1 0 99360 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_1080
timestamp 1
transform 1 0 100464 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_3
timestamp 1
transform 1 0 1380 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1056
timestamp 1636968456
transform 1 0 98256 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_1068
timestamp 1636968456
transform 1 0 99360 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_1080
timestamp 1
transform 1 0 100464 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_3
timestamp 1
transform 1 0 1380 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1056
timestamp 1636968456
transform 1 0 98256 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_1068
timestamp 1636968456
transform 1 0 99360 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_1080
timestamp 1
transform 1 0 100464 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_3
timestamp 1
transform 1 0 1380 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1056
timestamp 1636968456
transform 1 0 98256 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_1068
timestamp 1636968456
transform 1 0 99360 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_1080
timestamp 1
transform 1 0 100464 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_3
timestamp 1
transform 1 0 1380 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1056
timestamp 1636968456
transform 1 0 98256 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_1068
timestamp 1636968456
transform 1 0 99360 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_1080
timestamp 1
transform 1 0 100464 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_3
timestamp 1
transform 1 0 1380 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_1063
timestamp 1636968456
transform 1 0 98900 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_1075
timestamp 1
transform 1 0 100004 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_30_3
timestamp 1
transform 1 0 1380 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1056
timestamp 1636968456
transform 1 0 98256 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_1068
timestamp 1636968456
transform 1 0 99360 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_1080
timestamp 1
transform 1 0 100464 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_3
timestamp 1
transform 1 0 1380 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_1056
timestamp 1
transform 1 0 98256 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_1066
timestamp 1636968456
transform 1 0 99176 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_1078
timestamp 1
transform 1 0 100280 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_32_3
timestamp 1
transform 1 0 1380 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_1077
timestamp 1
transform 1 0 100188 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_33_3
timestamp 1
transform 1 0 1380 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1056
timestamp 1636968456
transform 1 0 98256 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_1068
timestamp 1636968456
transform 1 0 99360 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_1080
timestamp 1
transform 1 0 100464 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_34_3
timestamp 1
transform 1 0 1380 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1056
timestamp 1636968456
transform 1 0 98256 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_1068
timestamp 1636968456
transform 1 0 99360 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_1080
timestamp 1
transform 1 0 100464 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_3
timestamp 1
transform 1 0 1380 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1056
timestamp 1636968456
transform 1 0 98256 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_1068
timestamp 1636968456
transform 1 0 99360 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_1080
timestamp 1
transform 1 0 100464 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_36_3
timestamp 1
transform 1 0 1380 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_1061
timestamp 1636968456
transform 1 0 98716 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_1073
timestamp 1
transform 1 0 99820 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_3
timestamp 1
transform 1 0 1380 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_1065
timestamp 1
transform 1 0 99084 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_1070
timestamp 1
transform 1 0 99544 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_1078
timestamp 1
transform 1 0 100280 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_38_3
timestamp 1
transform 1 0 1380 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1056
timestamp 1636968456
transform 1 0 98256 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_1068
timestamp 1636968456
transform 1 0 99360 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_1080
timestamp 1
transform 1 0 100464 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_39_3
timestamp 1
transform 1 0 1380 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_1064
timestamp 1636968456
transform 1 0 98992 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_1076
timestamp 1
transform 1 0 100096 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_1080
timestamp 1
transform 1 0 100464 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_40_3
timestamp 1
transform 1 0 1380 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_40_1056
timestamp 1
transform 1 0 98256 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_1060
timestamp 1636968456
transform 1 0 98624 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_1072
timestamp 1
transform 1 0 99728 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_1080
timestamp 1
transform 1 0 100464 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_41_3
timestamp 1
transform 1 0 1380 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_41_1056
timestamp 1
transform 1 0 98256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_41_1078
timestamp 1
transform 1 0 100280 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_42_3
timestamp 1
transform 1 0 1380 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_1077
timestamp 1
transform 1 0 100188 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_43_3
timestamp 1
transform 1 0 1380 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_43_1056
timestamp 1
transform 1 0 98256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_1073
timestamp 1
transform 1 0 99820 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_3
timestamp 1
transform 1 0 1380 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_1056
timestamp 1
transform 1 0 98256 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_1064
timestamp 1636968456
transform 1 0 98992 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_1076
timestamp 1
transform 1 0 100096 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_45_3
timestamp 1
transform 1 0 1380 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1056
timestamp 1636968456
transform 1 0 98256 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_1068
timestamp 1636968456
transform 1 0 99360 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_1080
timestamp 1
transform 1 0 100464 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_46_3
timestamp 1
transform 1 0 1380 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_46_1056
timestamp 1
transform 1 0 98256 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_1064
timestamp 1
transform 1 0 98992 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_1075
timestamp 1
transform 1 0 100004 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_47_3
timestamp 1
transform 1 0 1380 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_1056
timestamp 1636968456
transform 1 0 98256 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_1068
timestamp 1636968456
transform 1 0 99360 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_1080
timestamp 1
transform 1 0 100464 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_48_3
timestamp 1
transform 1 0 1380 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_48_1056
timestamp 1636968456
transform 1 0 98256 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_1068
timestamp 1636968456
transform 1 0 99360 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_1080
timestamp 1
transform 1 0 100464 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_49_3
timestamp 1
transform 1 0 1380 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_49_1056
timestamp 1
transform 1 0 98256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_1060
timestamp 1
transform 1 0 98624 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_1077
timestamp 1
transform 1 0 100188 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_50_3
timestamp 1
transform 1 0 1380 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_1059
timestamp 1636968456
transform 1 0 98532 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_1071
timestamp 1
transform 1 0 99636 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_1079
timestamp 1
transform 1 0 100372 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_51_3
timestamp 1
transform 1 0 1380 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_1056
timestamp 1
transform 1 0 98256 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_1060
timestamp 1
transform 1 0 98624 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_1069
timestamp 1636968456
transform 1 0 99452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_3
timestamp 1
transform 1 0 1380 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_1076
timestamp 1
transform 1 0 100096 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_1080
timestamp 1
transform 1 0 100464 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_53_3
timestamp 1
transform 1 0 1380 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_1056
timestamp 1636968456
transform 1 0 98256 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_1068
timestamp 1636968456
transform 1 0 99360 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_1080
timestamp 1
transform 1 0 100464 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_54_3
timestamp 1
transform 1 0 1380 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_1077
timestamp 1
transform 1 0 100188 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_55_3
timestamp 1
transform 1 0 1380 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_55_1056
timestamp 1636968456
transform 1 0 98256 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_1068
timestamp 1636968456
transform 1 0 99360 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_1080
timestamp 1
transform 1 0 100464 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_56_3
timestamp 1
transform 1 0 1380 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_56_1056
timestamp 1636968456
transform 1 0 98256 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_1068
timestamp 1636968456
transform 1 0 99360 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_1080
timestamp 1
transform 1 0 100464 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_57_3
timestamp 1
transform 1 0 1380 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_1056
timestamp 1636968456
transform 1 0 98256 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_1068
timestamp 1636968456
transform 1 0 99360 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_1080
timestamp 1
transform 1 0 100464 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_58_3
timestamp 1
transform 1 0 1380 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_58_1056
timestamp 1636968456
transform 1 0 98256 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_1068
timestamp 1636968456
transform 1 0 99360 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_1080
timestamp 1
transform 1 0 100464 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_59_3
timestamp 1
transform 1 0 1380 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_59_1059
timestamp 1636968456
transform 1 0 98532 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_1071
timestamp 1
transform 1 0 99636 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_1079
timestamp 1
transform 1 0 100372 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_60_3
timestamp 1
transform 1 0 1380 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_60_1056
timestamp 1636968456
transform 1 0 98256 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_1068
timestamp 1636968456
transform 1 0 99360 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_1080
timestamp 1
transform 1 0 100464 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_61_3
timestamp 1
transform 1 0 1380 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_61_1059
timestamp 1636968456
transform 1 0 98532 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_1071
timestamp 1
transform 1 0 99636 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_1079
timestamp 1
transform 1 0 100372 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_62_3
timestamp 1
transform 1 0 1380 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_62_1056
timestamp 1636968456
transform 1 0 98256 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_1068
timestamp 1636968456
transform 1 0 99360 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_1080
timestamp 1
transform 1 0 100464 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_63_3
timestamp 1
transform 1 0 1380 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_63_1056
timestamp 1636968456
transform 1 0 98256 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_1068
timestamp 1636968456
transform 1 0 99360 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_1080
timestamp 1
transform 1 0 100464 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_64_3
timestamp 1
transform 1 0 1380 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_1056
timestamp 1636968456
transform 1 0 98256 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_1068
timestamp 1636968456
transform 1 0 99360 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_1080
timestamp 1
transform 1 0 100464 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_65_3
timestamp 1
transform 1 0 1380 0 -1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_65_1056
timestamp 1636968456
transform 1 0 98256 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_1068
timestamp 1636968456
transform 1 0 99360 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_1080
timestamp 1
transform 1 0 100464 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_66_3
timestamp 1
transform 1 0 1380 0 1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_66_1056
timestamp 1636968456
transform 1 0 98256 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_1068
timestamp 1636968456
transform 1 0 99360 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_1080
timestamp 1
transform 1 0 100464 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_67_3
timestamp 1
transform 1 0 1380 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_67_1056
timestamp 1636968456
transform 1 0 98256 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_1068
timestamp 1636968456
transform 1 0 99360 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_1080
timestamp 1
transform 1 0 100464 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_68_3
timestamp 1
transform 1 0 1380 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_68_1056
timestamp 1636968456
transform 1 0 98256 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_1068
timestamp 1636968456
transform 1 0 99360 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_1080
timestamp 1
transform 1 0 100464 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_69_3
timestamp 1
transform 1 0 1380 0 -1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_69_1056
timestamp 1636968456
transform 1 0 98256 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_1068
timestamp 1636968456
transform 1 0 99360 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_69_1080
timestamp 1
transform 1 0 100464 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_70_3
timestamp 1
transform 1 0 1380 0 1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_70_1059
timestamp 1636968456
transform 1 0 98532 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_1071
timestamp 1
transform 1 0 99636 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_70_1079
timestamp 1
transform 1 0 100372 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_71_3
timestamp 1
transform 1 0 1380 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_71_1077
timestamp 1
transform 1 0 100188 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_72_3
timestamp 1
transform 1 0 1380 0 1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_72_1056
timestamp 1636968456
transform 1 0 98256 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_1068
timestamp 1636968456
transform 1 0 99360 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_1080
timestamp 1
transform 1 0 100464 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_73_3
timestamp 1
transform 1 0 1380 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_73_1056
timestamp 1636968456
transform 1 0 98256 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_1068
timestamp 1636968456
transform 1 0 99360 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_73_1080
timestamp 1
transform 1 0 100464 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_74_3
timestamp 1
transform 1 0 1380 0 1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_74_1056
timestamp 1636968456
transform 1 0 98256 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_1068
timestamp 1636968456
transform 1 0 99360 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_1080
timestamp 1
transform 1 0 100464 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_75_3
timestamp 1
transform 1 0 1380 0 -1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_75_1059
timestamp 1636968456
transform 1 0 98532 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_1071
timestamp 1
transform 1 0 99636 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_75_1079
timestamp 1
transform 1 0 100372 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_76_3
timestamp 1
transform 1 0 1380 0 1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_76_1056
timestamp 1636968456
transform 1 0 98256 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_1068
timestamp 1636968456
transform 1 0 99360 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_1080
timestamp 1
transform 1 0 100464 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_77_3
timestamp 1
transform 1 0 1380 0 -1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_77_1056
timestamp 1636968456
transform 1 0 98256 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_1068
timestamp 1636968456
transform 1 0 99360 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_77_1080
timestamp 1
transform 1 0 100464 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_78_3
timestamp 1
transform 1 0 1380 0 1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_78_1062
timestamp 1636968456
transform 1 0 98808 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_1074
timestamp 1
transform 1 0 99912 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_1080
timestamp 1
transform 1 0 100464 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_79_3
timestamp 1
transform 1 0 1380 0 -1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_79_1056
timestamp 1636968456
transform 1 0 98256 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_1068
timestamp 1636968456
transform 1 0 99360 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_79_1080
timestamp 1
transform 1 0 100464 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_80_3
timestamp 1
transform 1 0 1380 0 1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_80_1060
timestamp 1636968456
transform 1 0 98624 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_1072
timestamp 1
transform 1 0 99728 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_1080
timestamp 1
transform 1 0 100464 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_81_3
timestamp 1
transform 1 0 1380 0 -1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_81_1056
timestamp 1636968456
transform 1 0 98256 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_1068
timestamp 1636968456
transform 1 0 99360 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_81_1080
timestamp 1
transform 1 0 100464 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_82_3
timestamp 1
transform 1 0 1380 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_82_1056
timestamp 1636968456
transform 1 0 98256 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_1068
timestamp 1636968456
transform 1 0 99360 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_1080
timestamp 1
transform 1 0 100464 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_83_3
timestamp 1
transform 1 0 1380 0 -1 47872
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_83_1056
timestamp 1636968456
transform 1 0 98256 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_1068
timestamp 1636968456
transform 1 0 99360 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_83_1080
timestamp 1
transform 1 0 100464 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_84_3
timestamp 1
transform 1 0 1380 0 1 47872
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_84_1056
timestamp 1636968456
transform 1 0 98256 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_1068
timestamp 1636968456
transform 1 0 99360 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_1080
timestamp 1
transform 1 0 100464 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_85_3
timestamp 1
transform 1 0 1380 0 -1 48960
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_85_1056
timestamp 1636968456
transform 1 0 98256 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_1068
timestamp 1636968456
transform 1 0 99360 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_85_1080
timestamp 1
transform 1 0 100464 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_86_3
timestamp 1
transform 1 0 1380 0 1 48960
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_86_1056
timestamp 1636968456
transform 1 0 98256 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_1068
timestamp 1636968456
transform 1 0 99360 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_1080
timestamp 1
transform 1 0 100464 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_87_3
timestamp 1
transform 1 0 1380 0 -1 50048
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_87_1056
timestamp 1636968456
transform 1 0 98256 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_1068
timestamp 1636968456
transform 1 0 99360 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_87_1080
timestamp 1
transform 1 0 100464 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_88_3
timestamp 1
transform 1 0 1380 0 1 50048
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_88_1056
timestamp 1636968456
transform 1 0 98256 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_1068
timestamp 1636968456
transform 1 0 99360 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_88_1080
timestamp 1
transform 1 0 100464 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_89_3
timestamp 1
transform 1 0 1380 0 -1 51136
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_89_1056
timestamp 1636968456
transform 1 0 98256 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_1068
timestamp 1636968456
transform 1 0 99360 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_89_1080
timestamp 1
transform 1 0 100464 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_90_3
timestamp 1
transform 1 0 1380 0 1 51136
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_90_1056
timestamp 1636968456
transform 1 0 98256 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_1068
timestamp 1636968456
transform 1 0 99360 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_90_1080
timestamp 1
transform 1 0 100464 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_91_3
timestamp 1
transform 1 0 1380 0 -1 52224
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_91_1056
timestamp 1636968456
transform 1 0 98256 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_1068
timestamp 1636968456
transform 1 0 99360 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_91_1080
timestamp 1
transform 1 0 100464 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_92_3
timestamp 1
transform 1 0 1380 0 1 52224
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_92_1056
timestamp 1636968456
transform 1 0 98256 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_1068
timestamp 1636968456
transform 1 0 99360 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_92_1080
timestamp 1
transform 1 0 100464 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_93_3
timestamp 1
transform 1 0 1380 0 -1 53312
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_93_1056
timestamp 1636968456
transform 1 0 98256 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_1068
timestamp 1636968456
transform 1 0 99360 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_93_1080
timestamp 1
transform 1 0 100464 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_94_3
timestamp 1
transform 1 0 1380 0 1 53312
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_94_1056
timestamp 1636968456
transform 1 0 98256 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_1068
timestamp 1636968456
transform 1 0 99360 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_94_1080
timestamp 1
transform 1 0 100464 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_95_3
timestamp 1
transform 1 0 1380 0 -1 54400
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_95_1059
timestamp 1636968456
transform 1 0 98532 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_95_1071
timestamp 1
transform 1 0 99636 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_95_1079
timestamp 1
transform 1 0 100372 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_96_3
timestamp 1
transform 1 0 1380 0 1 54400
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_96_1056
timestamp 1636968456
transform 1 0 98256 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_1068
timestamp 1636968456
transform 1 0 99360 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_96_1080
timestamp 1
transform 1 0 100464 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_97_3
timestamp 1
transform 1 0 1380 0 -1 55488
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_97_1056
timestamp 1636968456
transform 1 0 98256 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_1068
timestamp 1636968456
transform 1 0 99360 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_97_1080
timestamp 1
transform 1 0 100464 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_98_3
timestamp 1
transform 1 0 1380 0 1 55488
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_98_1056
timestamp 1636968456
transform 1 0 98256 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_1068
timestamp 1636968456
transform 1 0 99360 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_98_1080
timestamp 1
transform 1 0 100464 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_99_3
timestamp 1
transform 1 0 1380 0 -1 56576
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_99_1056
timestamp 1636968456
transform 1 0 98256 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_1068
timestamp 1636968456
transform 1 0 99360 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_99_1080
timestamp 1
transform 1 0 100464 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_100_3
timestamp 1
transform 1 0 1380 0 1 56576
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_100_1056
timestamp 1636968456
transform 1 0 98256 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_1068
timestamp 1636968456
transform 1 0 99360 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_100_1080
timestamp 1
transform 1 0 100464 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_101_3
timestamp 1
transform 1 0 1380 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_1056
timestamp 1636968456
transform 1 0 98256 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_1068
timestamp 1636968456
transform 1 0 99360 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_101_1080
timestamp 1
transform 1 0 100464 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_102_3
timestamp 1
transform 1 0 1380 0 1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_102_1056
timestamp 1636968456
transform 1 0 98256 0 1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_1068
timestamp 1636968456
transform 1 0 99360 0 1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_102_1080
timestamp 1
transform 1 0 100464 0 1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_103_3
timestamp 1
transform 1 0 1380 0 -1 58752
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_103_1056
timestamp 1636968456
transform 1 0 98256 0 -1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_1068
timestamp 1636968456
transform 1 0 99360 0 -1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_103_1080
timestamp 1
transform 1 0 100464 0 -1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_104_3
timestamp 1
transform 1 0 1380 0 1 58752
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_104_1056
timestamp 1636968456
transform 1 0 98256 0 1 58752
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_1068
timestamp 1636968456
transform 1 0 99360 0 1 58752
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_104_1080
timestamp 1
transform 1 0 100464 0 1 58752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_105_3
timestamp 1
transform 1 0 1380 0 -1 59840
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_105_1056
timestamp 1636968456
transform 1 0 98256 0 -1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_1068
timestamp 1636968456
transform 1 0 99360 0 -1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_105_1080
timestamp 1
transform 1 0 100464 0 -1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_3
timestamp 1636968456
transform 1 0 1380 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_15
timestamp 1636968456
transform 1 0 2484 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_106_27
timestamp 1
transform 1 0 3588 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_29
timestamp 1636968456
transform 1 0 3772 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_41
timestamp 1636968456
transform 1 0 4876 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_106_53
timestamp 1
transform 1 0 5980 0 1 59840
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_106_57
timestamp 1636968456
transform 1 0 6348 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_69
timestamp 1636968456
transform 1 0 7452 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_106_81
timestamp 1
transform 1 0 8556 0 1 59840
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_106_85
timestamp 1636968456
transform 1 0 8924 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_97
timestamp 1636968456
transform 1 0 10028 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_106_109
timestamp 1
transform 1 0 11132 0 1 59840
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_106_113
timestamp 1636968456
transform 1 0 11500 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_125
timestamp 1636968456
transform 1 0 12604 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_106_137
timestamp 1
transform 1 0 13708 0 1 59840
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_106_141
timestamp 1636968456
transform 1 0 14076 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_153
timestamp 1636968456
transform 1 0 15180 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_106_165
timestamp 1
transform 1 0 16284 0 1 59840
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_106_169
timestamp 1636968456
transform 1 0 16652 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_181
timestamp 1636968456
transform 1 0 17756 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_106_193
timestamp 1
transform 1 0 18860 0 1 59840
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_106_197
timestamp 1636968456
transform 1 0 19228 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_209
timestamp 1636968456
transform 1 0 20332 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_106_221
timestamp 1
transform 1 0 21436 0 1 59840
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_106_225
timestamp 1636968456
transform 1 0 21804 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_237
timestamp 1636968456
transform 1 0 22908 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_106_249
timestamp 1
transform 1 0 24012 0 1 59840
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_106_253
timestamp 1636968456
transform 1 0 24380 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_265
timestamp 1636968456
transform 1 0 25484 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_106_277
timestamp 1
transform 1 0 26588 0 1 59840
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_106_281
timestamp 1636968456
transform 1 0 26956 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_293
timestamp 1636968456
transform 1 0 28060 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_106_305
timestamp 1
transform 1 0 29164 0 1 59840
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_106_309
timestamp 1636968456
transform 1 0 29532 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_321
timestamp 1636968456
transform 1 0 30636 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_106_333
timestamp 1
transform 1 0 31740 0 1 59840
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_106_337
timestamp 1636968456
transform 1 0 32108 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_349
timestamp 1636968456
transform 1 0 33212 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_106_361
timestamp 1
transform 1 0 34316 0 1 59840
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_106_365
timestamp 1636968456
transform 1 0 34684 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_377
timestamp 1636968456
transform 1 0 35788 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_106_389
timestamp 1
transform 1 0 36892 0 1 59840
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_106_393
timestamp 1636968456
transform 1 0 37260 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_405
timestamp 1636968456
transform 1 0 38364 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_106_417
timestamp 1
transform 1 0 39468 0 1 59840
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_106_421
timestamp 1636968456
transform 1 0 39836 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_433
timestamp 1636968456
transform 1 0 40940 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_106_445
timestamp 1
transform 1 0 42044 0 1 59840
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_106_449
timestamp 1636968456
transform 1 0 42412 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_461
timestamp 1636968456
transform 1 0 43516 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_106_473
timestamp 1
transform 1 0 44620 0 1 59840
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_106_477
timestamp 1636968456
transform 1 0 44988 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_489
timestamp 1636968456
transform 1 0 46092 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_106_501
timestamp 1
transform 1 0 47196 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_106_505
timestamp 1
transform 1 0 47564 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_531
timestamp 1
transform 1 0 49956 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_533
timestamp 1636968456
transform 1 0 50140 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_545
timestamp 1636968456
transform 1 0 51244 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_106_557
timestamp 1
transform 1 0 52348 0 1 59840
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_106_561
timestamp 1636968456
transform 1 0 52716 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_573
timestamp 1636968456
transform 1 0 53820 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_106_585
timestamp 1
transform 1 0 54924 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_106_609
timestamp 1
transform 1 0 57132 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_615
timestamp 1
transform 1 0 57684 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_617
timestamp 1636968456
transform 1 0 57868 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_629
timestamp 1636968456
transform 1 0 58972 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_106_641
timestamp 1
transform 1 0 60076 0 1 59840
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_106_645
timestamp 1636968456
transform 1 0 60444 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_657
timestamp 1636968456
transform 1 0 61548 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_106_669
timestamp 1
transform 1 0 62652 0 1 59840
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_106_673
timestamp 1636968456
transform 1 0 63020 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_685
timestamp 1636968456
transform 1 0 64124 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_106_697
timestamp 1
transform 1 0 65228 0 1 59840
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_106_701
timestamp 1636968456
transform 1 0 65596 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_713
timestamp 1636968456
transform 1 0 66700 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_106_725
timestamp 1
transform 1 0 67804 0 1 59840
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_106_729
timestamp 1636968456
transform 1 0 68172 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_741
timestamp 1636968456
transform 1 0 69276 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_106_753
timestamp 1
transform 1 0 70380 0 1 59840
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_106_757
timestamp 1636968456
transform 1 0 70748 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_769
timestamp 1636968456
transform 1 0 71852 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_106_781
timestamp 1
transform 1 0 72956 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_106_785
timestamp 1
transform 1 0 73324 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_106_809
timestamp 1
transform 1 0 75532 0 1 59840
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_106_813
timestamp 1636968456
transform 1 0 75900 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_825
timestamp 1636968456
transform 1 0 77004 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_106_837
timestamp 1
transform 1 0 78108 0 1 59840
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_106_841
timestamp 1636968456
transform 1 0 78476 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_106_853
timestamp 1
transform 1 0 79580 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_106_862
timestamp 1
transform 1 0 80408 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_106_869
timestamp 1
transform 1 0 81052 0 1 59840
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_106_875
timestamp 1
transform 1 0 81604 0 1 59840
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_879
timestamp 1636968456
transform 1 0 81972 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_106_891
timestamp 1
transform 1 0 83076 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_106_895
timestamp 1
transform 1 0 83444 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_106_897
timestamp 1
transform 1 0 83628 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_106_908
timestamp 1
transform 1 0 84640 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_106_912
timestamp 1
transform 1 0 85008 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_106_925
timestamp 1
transform 1 0 86204 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_106_948
timestamp 1
transform 1 0 88320 0 1 59840
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_106_953
timestamp 1636968456
transform 1 0 88780 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_965
timestamp 1636968456
transform 1 0 89884 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_106_977
timestamp 1
transform 1 0 90988 0 1 59840
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_106_981
timestamp 1636968456
transform 1 0 91356 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_993
timestamp 1636968456
transform 1 0 92460 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_106_1005
timestamp 1
transform 1 0 93564 0 1 59840
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_106_1009
timestamp 1636968456
transform 1 0 93932 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_1021
timestamp 1636968456
transform 1 0 95036 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_106_1033
timestamp 1
transform 1 0 96140 0 1 59840
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_106_1037
timestamp 1636968456
transform 1 0 96508 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_1049
timestamp 1636968456
transform 1 0 97612 0 1 59840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_106_1061
timestamp 1
transform 1 0 98716 0 1 59840
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_106_1065
timestamp 1636968456
transform 1 0 99084 0 1 59840
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_3
timestamp 1636968456
transform 1 0 1380 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_15
timestamp 1636968456
transform 1 0 2484 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_27
timestamp 1636968456
transform 1 0 3588 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_39
timestamp 1636968456
transform 1 0 4692 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_107_51
timestamp 1
transform 1 0 5796 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_107_55
timestamp 1
transform 1 0 6164 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_57
timestamp 1636968456
transform 1 0 6348 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_69
timestamp 1636968456
transform 1 0 7452 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_81
timestamp 1636968456
transform 1 0 8556 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_93
timestamp 1636968456
transform 1 0 9660 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_105
timestamp 1
transform 1 0 10764 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_111
timestamp 1
transform 1 0 11316 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_113
timestamp 1636968456
transform 1 0 11500 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_125
timestamp 1636968456
transform 1 0 12604 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_137
timestamp 1636968456
transform 1 0 13708 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_149
timestamp 1636968456
transform 1 0 14812 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_161
timestamp 1
transform 1 0 15916 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_167
timestamp 1
transform 1 0 16468 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_169
timestamp 1636968456
transform 1 0 16652 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_181
timestamp 1636968456
transform 1 0 17756 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_193
timestamp 1636968456
transform 1 0 18860 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_205
timestamp 1636968456
transform 1 0 19964 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_217
timestamp 1
transform 1 0 21068 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_223
timestamp 1
transform 1 0 21620 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_107_225
timestamp 1
transform 1 0 21804 0 -1 60928
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_107_253
timestamp 1636968456
transform 1 0 24380 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_265
timestamp 1636968456
transform 1 0 25484 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_107_277
timestamp 1
transform 1 0 26588 0 -1 60928
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_107_281
timestamp 1636968456
transform 1 0 26956 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_293
timestamp 1
transform 1 0 28060 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_107_301
timestamp 1
transform 1 0 28796 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_107_307
timestamp 1
transform 1 0 29348 0 -1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_107_315
timestamp 1
transform 1 0 30084 0 -1 60928
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_107_320
timestamp 1636968456
transform 1 0 30544 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_107_332
timestamp 1
transform 1 0 31648 0 -1 60928
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_107_337
timestamp 1636968456
transform 1 0 32108 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_349
timestamp 1636968456
transform 1 0 33212 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_361
timestamp 1636968456
transform 1 0 34316 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_373
timestamp 1636968456
transform 1 0 35420 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_385
timestamp 1
transform 1 0 36524 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_391
timestamp 1
transform 1 0 37076 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_393
timestamp 1636968456
transform 1 0 37260 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_405
timestamp 1636968456
transform 1 0 38364 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_417
timestamp 1636968456
transform 1 0 39468 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_429
timestamp 1636968456
transform 1 0 40572 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_441
timestamp 1
transform 1 0 41676 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_447
timestamp 1
transform 1 0 42228 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_449
timestamp 1636968456
transform 1 0 42412 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_461
timestamp 1636968456
transform 1 0 43516 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_473
timestamp 1636968456
transform 1 0 44620 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_485
timestamp 1636968456
transform 1 0 45724 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_497
timestamp 1
transform 1 0 46828 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_503
timestamp 1
transform 1 0 47380 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_107_505
timestamp 1
transform 1 0 47564 0 -1 60928
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_107_522
timestamp 1636968456
transform 1 0 49128 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_534
timestamp 1636968456
transform 1 0 50232 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_546
timestamp 1636968456
transform 1 0 51336 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_107_558
timestamp 1
transform 1 0 52440 0 -1 60928
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_107_561
timestamp 1636968456
transform 1 0 52716 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_573
timestamp 1636968456
transform 1 0 53820 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_585
timestamp 1636968456
transform 1 0 54924 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_597
timestamp 1636968456
transform 1 0 56028 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_609
timestamp 1
transform 1 0 57132 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_615
timestamp 1
transform 1 0 57684 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_617
timestamp 1636968456
transform 1 0 57868 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_629
timestamp 1636968456
transform 1 0 58972 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_641
timestamp 1636968456
transform 1 0 60076 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_653
timestamp 1636968456
transform 1 0 61180 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_665
timestamp 1
transform 1 0 62284 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_671
timestamp 1
transform 1 0 62836 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_673
timestamp 1636968456
transform 1 0 63020 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_685
timestamp 1636968456
transform 1 0 64124 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_697
timestamp 1636968456
transform 1 0 65228 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_709
timestamp 1636968456
transform 1 0 66332 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_721
timestamp 1
transform 1 0 67436 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_727
timestamp 1
transform 1 0 67988 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_729
timestamp 1636968456
transform 1 0 68172 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_741
timestamp 1636968456
transform 1 0 69276 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_753
timestamp 1636968456
transform 1 0 70380 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_765
timestamp 1636968456
transform 1 0 71484 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_777
timestamp 1
transform 1 0 72588 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_783
timestamp 1
transform 1 0 73140 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_785
timestamp 1636968456
transform 1 0 73324 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_797
timestamp 1636968456
transform 1 0 74428 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_809
timestamp 1636968456
transform 1 0 75532 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_107_821
timestamp 1
transform 1 0 76636 0 -1 60928
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_107_828
timestamp 1636968456
transform 1 0 77280 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_107_844
timestamp 1
transform 1 0 78752 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_107_848
timestamp 1
transform 1 0 79120 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_107_897
timestamp 1
transform 1 0 83628 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_107_944
timestamp 1
transform 1 0 87952 0 -1 60928
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_107_953
timestamp 1636968456
transform 1 0 88780 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_965
timestamp 1636968456
transform 1 0 89884 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_977
timestamp 1636968456
transform 1 0 90988 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_989
timestamp 1636968456
transform 1 0 92092 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_1001
timestamp 1
transform 1 0 93196 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_1007
timestamp 1
transform 1 0 93748 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_1009
timestamp 1636968456
transform 1 0 93932 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_1021
timestamp 1636968456
transform 1 0 95036 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_1033
timestamp 1636968456
transform 1 0 96140 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_1045
timestamp 1636968456
transform 1 0 97244 0 -1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_107_1057
timestamp 1
transform 1 0 98348 0 -1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_1063
timestamp 1
transform 1 0 98900 0 -1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_1065
timestamp 1636968456
transform 1 0 99084 0 -1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_3
timestamp 1636968456
transform 1 0 1380 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_15
timestamp 1636968456
transform 1 0 2484 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_108_27
timestamp 1
transform 1 0 3588 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_29
timestamp 1636968456
transform 1 0 3772 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_41
timestamp 1636968456
transform 1 0 4876 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_53
timestamp 1636968456
transform 1 0 5980 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_65
timestamp 1636968456
transform 1 0 7084 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_77
timestamp 1
transform 1 0 8188 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_83
timestamp 1
transform 1 0 8740 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_85
timestamp 1636968456
transform 1 0 8924 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_97
timestamp 1636968456
transform 1 0 10028 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_109
timestamp 1636968456
transform 1 0 11132 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_121
timestamp 1636968456
transform 1 0 12236 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_133
timestamp 1
transform 1 0 13340 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_139
timestamp 1
transform 1 0 13892 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_141
timestamp 1636968456
transform 1 0 14076 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_153
timestamp 1636968456
transform 1 0 15180 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_165
timestamp 1636968456
transform 1 0 16284 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_177
timestamp 1636968456
transform 1 0 17388 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_189
timestamp 1
transform 1 0 18492 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_195
timestamp 1
transform 1 0 19044 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_197
timestamp 1636968456
transform 1 0 19228 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_108_209
timestamp 1
transform 1 0 20332 0 1 60928
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_108_237
timestamp 1636968456
transform 1 0 22908 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_108_249
timestamp 1
transform 1 0 24012 0 1 60928
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_108_253
timestamp 1636968456
transform 1 0 24380 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_265
timestamp 1636968456
transform 1 0 25484 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_277
timestamp 1636968456
transform 1 0 26588 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_289
timestamp 1636968456
transform 1 0 27692 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_301
timestamp 1
transform 1 0 28796 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_307
timestamp 1
transform 1 0 29348 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_309
timestamp 1636968456
transform 1 0 29532 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_321
timestamp 1636968456
transform 1 0 30636 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_333
timestamp 1636968456
transform 1 0 31740 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_345
timestamp 1636968456
transform 1 0 32844 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_357
timestamp 1
transform 1 0 33948 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_363
timestamp 1
transform 1 0 34500 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_365
timestamp 1636968456
transform 1 0 34684 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_377
timestamp 1636968456
transform 1 0 35788 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_389
timestamp 1636968456
transform 1 0 36892 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_401
timestamp 1636968456
transform 1 0 37996 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_413
timestamp 1
transform 1 0 39100 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_419
timestamp 1
transform 1 0 39652 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_421
timestamp 1636968456
transform 1 0 39836 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_433
timestamp 1636968456
transform 1 0 40940 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_445
timestamp 1636968456
transform 1 0 42044 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_457
timestamp 1636968456
transform 1 0 43148 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_469
timestamp 1
transform 1 0 44252 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_475
timestamp 1
transform 1 0 44804 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_477
timestamp 1636968456
transform 1 0 44988 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_489
timestamp 1636968456
transform 1 0 46092 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_501
timestamp 1636968456
transform 1 0 47196 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_513
timestamp 1636968456
transform 1 0 48300 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_525
timestamp 1
transform 1 0 49404 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_531
timestamp 1
transform 1 0 49956 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_533
timestamp 1636968456
transform 1 0 50140 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_545
timestamp 1636968456
transform 1 0 51244 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_557
timestamp 1636968456
transform 1 0 52348 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_569
timestamp 1636968456
transform 1 0 53452 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_581
timestamp 1
transform 1 0 54556 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_587
timestamp 1
transform 1 0 55108 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_589
timestamp 1636968456
transform 1 0 55292 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_601
timestamp 1636968456
transform 1 0 56396 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_613
timestamp 1636968456
transform 1 0 57500 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_625
timestamp 1636968456
transform 1 0 58604 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_637
timestamp 1
transform 1 0 59708 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_643
timestamp 1
transform 1 0 60260 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_645
timestamp 1636968456
transform 1 0 60444 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_657
timestamp 1636968456
transform 1 0 61548 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_669
timestamp 1636968456
transform 1 0 62652 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_681
timestamp 1636968456
transform 1 0 63756 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_693
timestamp 1
transform 1 0 64860 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_699
timestamp 1
transform 1 0 65412 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_701
timestamp 1636968456
transform 1 0 65596 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_713
timestamp 1636968456
transform 1 0 66700 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_725
timestamp 1636968456
transform 1 0 67804 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_737
timestamp 1636968456
transform 1 0 68908 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_749
timestamp 1
transform 1 0 70012 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_755
timestamp 1
transform 1 0 70564 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_757
timestamp 1636968456
transform 1 0 70748 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_769
timestamp 1636968456
transform 1 0 71852 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_781
timestamp 1636968456
transform 1 0 72956 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_793
timestamp 1636968456
transform 1 0 74060 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_805
timestamp 1
transform 1 0 75164 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_811
timestamp 1
transform 1 0 75716 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_108_813
timestamp 1
transform 1 0 75900 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_108_821
timestamp 1
transform 1 0 76636 0 1 60928
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_108_867
timestamp 1
transform 1 0 80868 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_108_869
timestamp 1
transform 1 0 81052 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_108_877
timestamp 1
transform 1 0 81788 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_903
timestamp 1636968456
transform 1 0 84180 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_108_915
timestamp 1
transform 1 0 85284 0 1 60928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_108_923
timestamp 1
transform 1 0 86020 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_925
timestamp 1636968456
transform 1 0 86204 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_937
timestamp 1636968456
transform 1 0 87308 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_949
timestamp 1636968456
transform 1 0 88412 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_961
timestamp 1636968456
transform 1 0 89516 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_973
timestamp 1
transform 1 0 90620 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_979
timestamp 1
transform 1 0 91172 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_981
timestamp 1636968456
transform 1 0 91356 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_993
timestamp 1636968456
transform 1 0 92460 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_1005
timestamp 1636968456
transform 1 0 93564 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_1017
timestamp 1636968456
transform 1 0 94668 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_108_1029
timestamp 1
transform 1 0 95772 0 1 60928
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_108_1035
timestamp 1
transform 1 0 96324 0 1 60928
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_1037
timestamp 1636968456
transform 1 0 96508 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_1049
timestamp 1636968456
transform 1 0 97612 0 1 60928
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_1061
timestamp 1636968456
transform 1 0 98716 0 1 60928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_108_1073
timestamp 1
transform 1 0 99820 0 1 60928
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_109_7
timestamp 1636968456
transform 1 0 1748 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_19
timestamp 1636968456
transform 1 0 2852 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_31
timestamp 1636968456
transform 1 0 3956 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_43
timestamp 1636968456
transform 1 0 5060 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_109_55
timestamp 1
transform 1 0 6164 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_57
timestamp 1636968456
transform 1 0 6348 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_69
timestamp 1636968456
transform 1 0 7452 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_81
timestamp 1636968456
transform 1 0 8556 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_93
timestamp 1636968456
transform 1 0 9660 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_105
timestamp 1
transform 1 0 10764 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_111
timestamp 1
transform 1 0 11316 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_113
timestamp 1636968456
transform 1 0 11500 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_125
timestamp 1636968456
transform 1 0 12604 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_137
timestamp 1636968456
transform 1 0 13708 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_149
timestamp 1636968456
transform 1 0 14812 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_161
timestamp 1
transform 1 0 15916 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_167
timestamp 1
transform 1 0 16468 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_169
timestamp 1636968456
transform 1 0 16652 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_181
timestamp 1636968456
transform 1 0 17756 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_193
timestamp 1636968456
transform 1 0 18860 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_205
timestamp 1636968456
transform 1 0 19964 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_217
timestamp 1
transform 1 0 21068 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_223
timestamp 1
transform 1 0 21620 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_225
timestamp 1636968456
transform 1 0 21804 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_237
timestamp 1636968456
transform 1 0 22908 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_249
timestamp 1636968456
transform 1 0 24012 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_261
timestamp 1636968456
transform 1 0 25116 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_273
timestamp 1
transform 1 0 26220 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_279
timestamp 1
transform 1 0 26772 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_281
timestamp 1636968456
transform 1 0 26956 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_293
timestamp 1636968456
transform 1 0 28060 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_305
timestamp 1636968456
transform 1 0 29164 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_317
timestamp 1636968456
transform 1 0 30268 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_329
timestamp 1
transform 1 0 31372 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_335
timestamp 1
transform 1 0 31924 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_337
timestamp 1636968456
transform 1 0 32108 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_349
timestamp 1636968456
transform 1 0 33212 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_361
timestamp 1636968456
transform 1 0 34316 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_373
timestamp 1636968456
transform 1 0 35420 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_385
timestamp 1
transform 1 0 36524 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_391
timestamp 1
transform 1 0 37076 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_393
timestamp 1636968456
transform 1 0 37260 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_405
timestamp 1636968456
transform 1 0 38364 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_417
timestamp 1636968456
transform 1 0 39468 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_429
timestamp 1636968456
transform 1 0 40572 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_441
timestamp 1
transform 1 0 41676 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_447
timestamp 1
transform 1 0 42228 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_449
timestamp 1636968456
transform 1 0 42412 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_461
timestamp 1636968456
transform 1 0 43516 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_473
timestamp 1636968456
transform 1 0 44620 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_485
timestamp 1636968456
transform 1 0 45724 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_497
timestamp 1
transform 1 0 46828 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_503
timestamp 1
transform 1 0 47380 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_505
timestamp 1636968456
transform 1 0 47564 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_517
timestamp 1636968456
transform 1 0 48668 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_529
timestamp 1636968456
transform 1 0 49772 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_541
timestamp 1636968456
transform 1 0 50876 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_553
timestamp 1
transform 1 0 51980 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_559
timestamp 1
transform 1 0 52532 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_561
timestamp 1636968456
transform 1 0 52716 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_573
timestamp 1636968456
transform 1 0 53820 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_585
timestamp 1636968456
transform 1 0 54924 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_597
timestamp 1636968456
transform 1 0 56028 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_609
timestamp 1
transform 1 0 57132 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_615
timestamp 1
transform 1 0 57684 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_617
timestamp 1636968456
transform 1 0 57868 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_629
timestamp 1636968456
transform 1 0 58972 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_641
timestamp 1636968456
transform 1 0 60076 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_653
timestamp 1636968456
transform 1 0 61180 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_665
timestamp 1
transform 1 0 62284 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_671
timestamp 1
transform 1 0 62836 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_673
timestamp 1636968456
transform 1 0 63020 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_685
timestamp 1636968456
transform 1 0 64124 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_697
timestamp 1636968456
transform 1 0 65228 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_709
timestamp 1636968456
transform 1 0 66332 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_721
timestamp 1
transform 1 0 67436 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_727
timestamp 1
transform 1 0 67988 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_729
timestamp 1636968456
transform 1 0 68172 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_741
timestamp 1636968456
transform 1 0 69276 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_753
timestamp 1636968456
transform 1 0 70380 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_765
timestamp 1636968456
transform 1 0 71484 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_777
timestamp 1
transform 1 0 72588 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_783
timestamp 1
transform 1 0 73140 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_785
timestamp 1636968456
transform 1 0 73324 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_797
timestamp 1636968456
transform 1 0 74428 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_809
timestamp 1636968456
transform 1 0 75532 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_821
timestamp 1636968456
transform 1 0 76636 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_833
timestamp 1
transform 1 0 77740 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_839
timestamp 1
transform 1 0 78292 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_841
timestamp 1636968456
transform 1 0 78476 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_853
timestamp 1636968456
transform 1 0 79580 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_865
timestamp 1636968456
transform 1 0 80684 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_877
timestamp 1636968456
transform 1 0 81788 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_889
timestamp 1
transform 1 0 82892 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_895
timestamp 1
transform 1 0 83444 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_897
timestamp 1636968456
transform 1 0 83628 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_909
timestamp 1636968456
transform 1 0 84732 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_921
timestamp 1636968456
transform 1 0 85836 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_933
timestamp 1636968456
transform 1 0 86940 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_945
timestamp 1
transform 1 0 88044 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_951
timestamp 1
transform 1 0 88596 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_953
timestamp 1636968456
transform 1 0 88780 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_965
timestamp 1636968456
transform 1 0 89884 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_977
timestamp 1636968456
transform 1 0 90988 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_989
timestamp 1636968456
transform 1 0 92092 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_1001
timestamp 1
transform 1 0 93196 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_1007
timestamp 1
transform 1 0 93748 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_1009
timestamp 1636968456
transform 1 0 93932 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_1021
timestamp 1636968456
transform 1 0 95036 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_1033
timestamp 1636968456
transform 1 0 96140 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_1045
timestamp 1636968456
transform 1 0 97244 0 -1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_1057
timestamp 1
transform 1 0 98348 0 -1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_109_1063
timestamp 1
transform 1 0 98900 0 -1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_1065
timestamp 1636968456
transform 1 0 99084 0 -1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_9
timestamp 1636968456
transform 1 0 1932 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_21
timestamp 1
transform 1 0 3036 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_27
timestamp 1
transform 1 0 3588 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_29
timestamp 1636968456
transform 1 0 3772 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_41
timestamp 1636968456
transform 1 0 4876 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_53
timestamp 1636968456
transform 1 0 5980 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_65
timestamp 1636968456
transform 1 0 7084 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_77
timestamp 1
transform 1 0 8188 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_83
timestamp 1
transform 1 0 8740 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_85
timestamp 1636968456
transform 1 0 8924 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_97
timestamp 1636968456
transform 1 0 10028 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_109
timestamp 1636968456
transform 1 0 11132 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_121
timestamp 1636968456
transform 1 0 12236 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_133
timestamp 1
transform 1 0 13340 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_139
timestamp 1
transform 1 0 13892 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_141
timestamp 1636968456
transform 1 0 14076 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_153
timestamp 1636968456
transform 1 0 15180 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_165
timestamp 1636968456
transform 1 0 16284 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_177
timestamp 1636968456
transform 1 0 17388 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_189
timestamp 1
transform 1 0 18492 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_195
timestamp 1
transform 1 0 19044 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_197
timestamp 1636968456
transform 1 0 19228 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_209
timestamp 1636968456
transform 1 0 20332 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_221
timestamp 1636968456
transform 1 0 21436 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_233
timestamp 1636968456
transform 1 0 22540 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_245
timestamp 1
transform 1 0 23644 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_251
timestamp 1
transform 1 0 24196 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_253
timestamp 1636968456
transform 1 0 24380 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_265
timestamp 1636968456
transform 1 0 25484 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_277
timestamp 1636968456
transform 1 0 26588 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_289
timestamp 1636968456
transform 1 0 27692 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_301
timestamp 1
transform 1 0 28796 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_307
timestamp 1
transform 1 0 29348 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_309
timestamp 1636968456
transform 1 0 29532 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_321
timestamp 1636968456
transform 1 0 30636 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_333
timestamp 1636968456
transform 1 0 31740 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_345
timestamp 1636968456
transform 1 0 32844 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_357
timestamp 1
transform 1 0 33948 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_363
timestamp 1
transform 1 0 34500 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_365
timestamp 1636968456
transform 1 0 34684 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_377
timestamp 1636968456
transform 1 0 35788 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_389
timestamp 1636968456
transform 1 0 36892 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_401
timestamp 1636968456
transform 1 0 37996 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_413
timestamp 1
transform 1 0 39100 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_419
timestamp 1
transform 1 0 39652 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_421
timestamp 1636968456
transform 1 0 39836 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_433
timestamp 1636968456
transform 1 0 40940 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_445
timestamp 1636968456
transform 1 0 42044 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_457
timestamp 1636968456
transform 1 0 43148 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_469
timestamp 1
transform 1 0 44252 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_475
timestamp 1
transform 1 0 44804 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_477
timestamp 1636968456
transform 1 0 44988 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_489
timestamp 1636968456
transform 1 0 46092 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_501
timestamp 1636968456
transform 1 0 47196 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_513
timestamp 1636968456
transform 1 0 48300 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_525
timestamp 1
transform 1 0 49404 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_531
timestamp 1
transform 1 0 49956 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_533
timestamp 1636968456
transform 1 0 50140 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_545
timestamp 1636968456
transform 1 0 51244 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_557
timestamp 1636968456
transform 1 0 52348 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_569
timestamp 1636968456
transform 1 0 53452 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_581
timestamp 1
transform 1 0 54556 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_587
timestamp 1
transform 1 0 55108 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_589
timestamp 1636968456
transform 1 0 55292 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_601
timestamp 1636968456
transform 1 0 56396 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_613
timestamp 1636968456
transform 1 0 57500 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_625
timestamp 1636968456
transform 1 0 58604 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_637
timestamp 1
transform 1 0 59708 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_643
timestamp 1
transform 1 0 60260 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_645
timestamp 1636968456
transform 1 0 60444 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_657
timestamp 1636968456
transform 1 0 61548 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_669
timestamp 1636968456
transform 1 0 62652 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_681
timestamp 1636968456
transform 1 0 63756 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_693
timestamp 1
transform 1 0 64860 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_699
timestamp 1
transform 1 0 65412 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_701
timestamp 1636968456
transform 1 0 65596 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_713
timestamp 1636968456
transform 1 0 66700 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_725
timestamp 1636968456
transform 1 0 67804 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_737
timestamp 1636968456
transform 1 0 68908 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_749
timestamp 1
transform 1 0 70012 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_755
timestamp 1
transform 1 0 70564 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_757
timestamp 1636968456
transform 1 0 70748 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_769
timestamp 1636968456
transform 1 0 71852 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_781
timestamp 1636968456
transform 1 0 72956 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_793
timestamp 1636968456
transform 1 0 74060 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_805
timestamp 1
transform 1 0 75164 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_811
timestamp 1
transform 1 0 75716 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_813
timestamp 1636968456
transform 1 0 75900 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_825
timestamp 1636968456
transform 1 0 77004 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_837
timestamp 1636968456
transform 1 0 78108 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_849
timestamp 1636968456
transform 1 0 79212 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_861
timestamp 1
transform 1 0 80316 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_867
timestamp 1
transform 1 0 80868 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_869
timestamp 1636968456
transform 1 0 81052 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_881
timestamp 1636968456
transform 1 0 82156 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_893
timestamp 1636968456
transform 1 0 83260 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_905
timestamp 1636968456
transform 1 0 84364 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_917
timestamp 1
transform 1 0 85468 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_923
timestamp 1
transform 1 0 86020 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_925
timestamp 1636968456
transform 1 0 86204 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_937
timestamp 1636968456
transform 1 0 87308 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_949
timestamp 1636968456
transform 1 0 88412 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_961
timestamp 1636968456
transform 1 0 89516 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_973
timestamp 1
transform 1 0 90620 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_979
timestamp 1
transform 1 0 91172 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_981
timestamp 1636968456
transform 1 0 91356 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_993
timestamp 1636968456
transform 1 0 92460 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_1005
timestamp 1636968456
transform 1 0 93564 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_1017
timestamp 1636968456
transform 1 0 94668 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_110_1029
timestamp 1
transform 1 0 95772 0 1 62016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_110_1035
timestamp 1
transform 1 0 96324 0 1 62016
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_1037
timestamp 1636968456
transform 1 0 96508 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_1049
timestamp 1636968456
transform 1 0 97612 0 1 62016
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_110_1061
timestamp 1636968456
transform 1 0 98716 0 1 62016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_110_1073
timestamp 1
transform 1 0 99820 0 1 62016
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_111_3
timestamp 1636968456
transform 1 0 1380 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_15
timestamp 1636968456
transform 1 0 2484 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_27
timestamp 1636968456
transform 1 0 3588 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_39
timestamp 1636968456
transform 1 0 4692 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_111_51
timestamp 1
transform 1 0 5796 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_111_55
timestamp 1
transform 1 0 6164 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_111_57
timestamp 1636968456
transform 1 0 6348 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_69
timestamp 1636968456
transform 1 0 7452 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_81
timestamp 1636968456
transform 1 0 8556 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_93
timestamp 1636968456
transform 1 0 9660 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_105
timestamp 1
transform 1 0 10764 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_111
timestamp 1
transform 1 0 11316 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_111_113
timestamp 1636968456
transform 1 0 11500 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_125
timestamp 1636968456
transform 1 0 12604 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_137
timestamp 1636968456
transform 1 0 13708 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_149
timestamp 1636968456
transform 1 0 14812 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_161
timestamp 1
transform 1 0 15916 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_167
timestamp 1
transform 1 0 16468 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_111_169
timestamp 1636968456
transform 1 0 16652 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_181
timestamp 1636968456
transform 1 0 17756 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_193
timestamp 1636968456
transform 1 0 18860 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_205
timestamp 1636968456
transform 1 0 19964 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_217
timestamp 1
transform 1 0 21068 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_223
timestamp 1
transform 1 0 21620 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_111_225
timestamp 1636968456
transform 1 0 21804 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_237
timestamp 1636968456
transform 1 0 22908 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_249
timestamp 1636968456
transform 1 0 24012 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_261
timestamp 1636968456
transform 1 0 25116 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_273
timestamp 1
transform 1 0 26220 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_279
timestamp 1
transform 1 0 26772 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_111_281
timestamp 1636968456
transform 1 0 26956 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_293
timestamp 1636968456
transform 1 0 28060 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_305
timestamp 1636968456
transform 1 0 29164 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_317
timestamp 1636968456
transform 1 0 30268 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_329
timestamp 1
transform 1 0 31372 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_335
timestamp 1
transform 1 0 31924 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_111_337
timestamp 1636968456
transform 1 0 32108 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_349
timestamp 1636968456
transform 1 0 33212 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_361
timestamp 1636968456
transform 1 0 34316 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_373
timestamp 1636968456
transform 1 0 35420 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_385
timestamp 1
transform 1 0 36524 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_391
timestamp 1
transform 1 0 37076 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_111_393
timestamp 1636968456
transform 1 0 37260 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_405
timestamp 1636968456
transform 1 0 38364 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_417
timestamp 1636968456
transform 1 0 39468 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_429
timestamp 1636968456
transform 1 0 40572 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_441
timestamp 1
transform 1 0 41676 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_447
timestamp 1
transform 1 0 42228 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_111_449
timestamp 1636968456
transform 1 0 42412 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_461
timestamp 1636968456
transform 1 0 43516 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_473
timestamp 1636968456
transform 1 0 44620 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_485
timestamp 1636968456
transform 1 0 45724 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_497
timestamp 1
transform 1 0 46828 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_503
timestamp 1
transform 1 0 47380 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_111_505
timestamp 1636968456
transform 1 0 47564 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_517
timestamp 1636968456
transform 1 0 48668 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_529
timestamp 1636968456
transform 1 0 49772 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_541
timestamp 1636968456
transform 1 0 50876 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_553
timestamp 1
transform 1 0 51980 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_559
timestamp 1
transform 1 0 52532 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_111_561
timestamp 1636968456
transform 1 0 52716 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_573
timestamp 1636968456
transform 1 0 53820 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_585
timestamp 1636968456
transform 1 0 54924 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_597
timestamp 1636968456
transform 1 0 56028 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_609
timestamp 1
transform 1 0 57132 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_615
timestamp 1
transform 1 0 57684 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_111_617
timestamp 1636968456
transform 1 0 57868 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_629
timestamp 1636968456
transform 1 0 58972 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_641
timestamp 1636968456
transform 1 0 60076 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_653
timestamp 1636968456
transform 1 0 61180 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_665
timestamp 1
transform 1 0 62284 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_671
timestamp 1
transform 1 0 62836 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_111_673
timestamp 1636968456
transform 1 0 63020 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_685
timestamp 1636968456
transform 1 0 64124 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_697
timestamp 1636968456
transform 1 0 65228 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_709
timestamp 1636968456
transform 1 0 66332 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_721
timestamp 1
transform 1 0 67436 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_727
timestamp 1
transform 1 0 67988 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_111_729
timestamp 1636968456
transform 1 0 68172 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_741
timestamp 1636968456
transform 1 0 69276 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_753
timestamp 1636968456
transform 1 0 70380 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_765
timestamp 1636968456
transform 1 0 71484 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_777
timestamp 1
transform 1 0 72588 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_783
timestamp 1
transform 1 0 73140 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_111_785
timestamp 1636968456
transform 1 0 73324 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_797
timestamp 1636968456
transform 1 0 74428 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_809
timestamp 1636968456
transform 1 0 75532 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_821
timestamp 1636968456
transform 1 0 76636 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_833
timestamp 1
transform 1 0 77740 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_839
timestamp 1
transform 1 0 78292 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_111_841
timestamp 1636968456
transform 1 0 78476 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_853
timestamp 1636968456
transform 1 0 79580 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_865
timestamp 1636968456
transform 1 0 80684 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_877
timestamp 1636968456
transform 1 0 81788 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_889
timestamp 1
transform 1 0 82892 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_895
timestamp 1
transform 1 0 83444 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_111_897
timestamp 1636968456
transform 1 0 83628 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_909
timestamp 1636968456
transform 1 0 84732 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_921
timestamp 1636968456
transform 1 0 85836 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_933
timestamp 1636968456
transform 1 0 86940 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_945
timestamp 1
transform 1 0 88044 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_951
timestamp 1
transform 1 0 88596 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_111_953
timestamp 1636968456
transform 1 0 88780 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_965
timestamp 1636968456
transform 1 0 89884 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_977
timestamp 1636968456
transform 1 0 90988 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_989
timestamp 1636968456
transform 1 0 92092 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_1001
timestamp 1
transform 1 0 93196 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_1007
timestamp 1
transform 1 0 93748 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_111_1009
timestamp 1636968456
transform 1 0 93932 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_1021
timestamp 1636968456
transform 1 0 95036 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_1033
timestamp 1636968456
transform 1 0 96140 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_1045
timestamp 1636968456
transform 1 0 97244 0 -1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_1057
timestamp 1
transform 1 0 98348 0 -1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_111_1063
timestamp 1
transform 1 0 98900 0 -1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_111_1065
timestamp 1636968456
transform 1 0 99084 0 -1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_3
timestamp 1636968456
transform 1 0 1380 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_15
timestamp 1636968456
transform 1 0 2484 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_112_27
timestamp 1
transform 1 0 3588 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_29
timestamp 1636968456
transform 1 0 3772 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_41
timestamp 1636968456
transform 1 0 4876 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_53
timestamp 1636968456
transform 1 0 5980 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_65
timestamp 1636968456
transform 1 0 7084 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_77
timestamp 1
transform 1 0 8188 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_83
timestamp 1
transform 1 0 8740 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_85
timestamp 1636968456
transform 1 0 8924 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_97
timestamp 1636968456
transform 1 0 10028 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_109
timestamp 1636968456
transform 1 0 11132 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_121
timestamp 1636968456
transform 1 0 12236 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_133
timestamp 1
transform 1 0 13340 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_139
timestamp 1
transform 1 0 13892 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_141
timestamp 1636968456
transform 1 0 14076 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_153
timestamp 1636968456
transform 1 0 15180 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_165
timestamp 1636968456
transform 1 0 16284 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_177
timestamp 1636968456
transform 1 0 17388 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_189
timestamp 1
transform 1 0 18492 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_195
timestamp 1
transform 1 0 19044 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_197
timestamp 1636968456
transform 1 0 19228 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_209
timestamp 1636968456
transform 1 0 20332 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_221
timestamp 1636968456
transform 1 0 21436 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_233
timestamp 1636968456
transform 1 0 22540 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_245
timestamp 1
transform 1 0 23644 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_251
timestamp 1
transform 1 0 24196 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_253
timestamp 1636968456
transform 1 0 24380 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_265
timestamp 1636968456
transform 1 0 25484 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_277
timestamp 1636968456
transform 1 0 26588 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_289
timestamp 1636968456
transform 1 0 27692 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_301
timestamp 1
transform 1 0 28796 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_307
timestamp 1
transform 1 0 29348 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_309
timestamp 1636968456
transform 1 0 29532 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_321
timestamp 1636968456
transform 1 0 30636 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_333
timestamp 1636968456
transform 1 0 31740 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_345
timestamp 1636968456
transform 1 0 32844 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_357
timestamp 1
transform 1 0 33948 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_363
timestamp 1
transform 1 0 34500 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_365
timestamp 1636968456
transform 1 0 34684 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_377
timestamp 1636968456
transform 1 0 35788 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_389
timestamp 1636968456
transform 1 0 36892 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_401
timestamp 1636968456
transform 1 0 37996 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_413
timestamp 1
transform 1 0 39100 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_419
timestamp 1
transform 1 0 39652 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_421
timestamp 1636968456
transform 1 0 39836 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_433
timestamp 1636968456
transform 1 0 40940 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_445
timestamp 1636968456
transform 1 0 42044 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_457
timestamp 1636968456
transform 1 0 43148 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_469
timestamp 1
transform 1 0 44252 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_475
timestamp 1
transform 1 0 44804 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_477
timestamp 1636968456
transform 1 0 44988 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_489
timestamp 1636968456
transform 1 0 46092 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_501
timestamp 1636968456
transform 1 0 47196 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_513
timestamp 1636968456
transform 1 0 48300 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_525
timestamp 1
transform 1 0 49404 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_531
timestamp 1
transform 1 0 49956 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_533
timestamp 1636968456
transform 1 0 50140 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_545
timestamp 1636968456
transform 1 0 51244 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_557
timestamp 1636968456
transform 1 0 52348 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_569
timestamp 1636968456
transform 1 0 53452 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_581
timestamp 1
transform 1 0 54556 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_587
timestamp 1
transform 1 0 55108 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_589
timestamp 1636968456
transform 1 0 55292 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_601
timestamp 1636968456
transform 1 0 56396 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_613
timestamp 1636968456
transform 1 0 57500 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_625
timestamp 1636968456
transform 1 0 58604 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_637
timestamp 1
transform 1 0 59708 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_643
timestamp 1
transform 1 0 60260 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_645
timestamp 1636968456
transform 1 0 60444 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_657
timestamp 1636968456
transform 1 0 61548 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_669
timestamp 1636968456
transform 1 0 62652 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_681
timestamp 1636968456
transform 1 0 63756 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_693
timestamp 1
transform 1 0 64860 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_699
timestamp 1
transform 1 0 65412 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_701
timestamp 1636968456
transform 1 0 65596 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_713
timestamp 1636968456
transform 1 0 66700 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_725
timestamp 1636968456
transform 1 0 67804 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_737
timestamp 1636968456
transform 1 0 68908 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_749
timestamp 1
transform 1 0 70012 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_755
timestamp 1
transform 1 0 70564 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_757
timestamp 1636968456
transform 1 0 70748 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_769
timestamp 1636968456
transform 1 0 71852 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_781
timestamp 1636968456
transform 1 0 72956 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_793
timestamp 1636968456
transform 1 0 74060 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_805
timestamp 1
transform 1 0 75164 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_811
timestamp 1
transform 1 0 75716 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_813
timestamp 1636968456
transform 1 0 75900 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_825
timestamp 1636968456
transform 1 0 77004 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_837
timestamp 1636968456
transform 1 0 78108 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_849
timestamp 1636968456
transform 1 0 79212 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_861
timestamp 1
transform 1 0 80316 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_867
timestamp 1
transform 1 0 80868 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_869
timestamp 1636968456
transform 1 0 81052 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_881
timestamp 1636968456
transform 1 0 82156 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_893
timestamp 1636968456
transform 1 0 83260 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_905
timestamp 1636968456
transform 1 0 84364 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_917
timestamp 1
transform 1 0 85468 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_923
timestamp 1
transform 1 0 86020 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_925
timestamp 1636968456
transform 1 0 86204 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_937
timestamp 1636968456
transform 1 0 87308 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_949
timestamp 1636968456
transform 1 0 88412 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_961
timestamp 1636968456
transform 1 0 89516 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_973
timestamp 1
transform 1 0 90620 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_979
timestamp 1
transform 1 0 91172 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_981
timestamp 1636968456
transform 1 0 91356 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_993
timestamp 1636968456
transform 1 0 92460 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_1005
timestamp 1636968456
transform 1 0 93564 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_1017
timestamp 1636968456
transform 1 0 94668 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_112_1029
timestamp 1
transform 1 0 95772 0 1 63104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_112_1035
timestamp 1
transform 1 0 96324 0 1 63104
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_1037
timestamp 1636968456
transform 1 0 96508 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_1049
timestamp 1636968456
transform 1 0 97612 0 1 63104
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_1061
timestamp 1636968456
transform 1 0 98716 0 1 63104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_112_1073
timestamp 1
transform 1 0 99820 0 1 63104
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_113_3
timestamp 1636968456
transform 1 0 1380 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_15
timestamp 1636968456
transform 1 0 2484 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_27
timestamp 1636968456
transform 1 0 3588 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_39
timestamp 1636968456
transform 1 0 4692 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_113_51
timestamp 1
transform 1 0 5796 0 -1 64192
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_113_55
timestamp 1
transform 1 0 6164 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_57
timestamp 1636968456
transform 1 0 6348 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_69
timestamp 1636968456
transform 1 0 7452 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_81
timestamp 1636968456
transform 1 0 8556 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_93
timestamp 1636968456
transform 1 0 9660 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_105
timestamp 1
transform 1 0 10764 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_111
timestamp 1
transform 1 0 11316 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_113
timestamp 1636968456
transform 1 0 11500 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_125
timestamp 1636968456
transform 1 0 12604 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_137
timestamp 1636968456
transform 1 0 13708 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_149
timestamp 1636968456
transform 1 0 14812 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_161
timestamp 1
transform 1 0 15916 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_167
timestamp 1
transform 1 0 16468 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_169
timestamp 1636968456
transform 1 0 16652 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_181
timestamp 1636968456
transform 1 0 17756 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_193
timestamp 1636968456
transform 1 0 18860 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_205
timestamp 1636968456
transform 1 0 19964 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_217
timestamp 1
transform 1 0 21068 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_223
timestamp 1
transform 1 0 21620 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_225
timestamp 1636968456
transform 1 0 21804 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_237
timestamp 1636968456
transform 1 0 22908 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_249
timestamp 1636968456
transform 1 0 24012 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_261
timestamp 1636968456
transform 1 0 25116 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_273
timestamp 1
transform 1 0 26220 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_279
timestamp 1
transform 1 0 26772 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_281
timestamp 1636968456
transform 1 0 26956 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_293
timestamp 1636968456
transform 1 0 28060 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_305
timestamp 1636968456
transform 1 0 29164 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_317
timestamp 1636968456
transform 1 0 30268 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_329
timestamp 1
transform 1 0 31372 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_335
timestamp 1
transform 1 0 31924 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_337
timestamp 1636968456
transform 1 0 32108 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_349
timestamp 1636968456
transform 1 0 33212 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_361
timestamp 1636968456
transform 1 0 34316 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_373
timestamp 1636968456
transform 1 0 35420 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_385
timestamp 1
transform 1 0 36524 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_391
timestamp 1
transform 1 0 37076 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_393
timestamp 1636968456
transform 1 0 37260 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_405
timestamp 1636968456
transform 1 0 38364 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_417
timestamp 1636968456
transform 1 0 39468 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_429
timestamp 1636968456
transform 1 0 40572 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_441
timestamp 1
transform 1 0 41676 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_447
timestamp 1
transform 1 0 42228 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_449
timestamp 1636968456
transform 1 0 42412 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_461
timestamp 1636968456
transform 1 0 43516 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_473
timestamp 1636968456
transform 1 0 44620 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_485
timestamp 1636968456
transform 1 0 45724 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_497
timestamp 1
transform 1 0 46828 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_503
timestamp 1
transform 1 0 47380 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_505
timestamp 1636968456
transform 1 0 47564 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_517
timestamp 1636968456
transform 1 0 48668 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_529
timestamp 1636968456
transform 1 0 49772 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_541
timestamp 1636968456
transform 1 0 50876 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_553
timestamp 1
transform 1 0 51980 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_559
timestamp 1
transform 1 0 52532 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_561
timestamp 1636968456
transform 1 0 52716 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_573
timestamp 1636968456
transform 1 0 53820 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_585
timestamp 1636968456
transform 1 0 54924 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_597
timestamp 1636968456
transform 1 0 56028 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_609
timestamp 1
transform 1 0 57132 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_615
timestamp 1
transform 1 0 57684 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_617
timestamp 1636968456
transform 1 0 57868 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_629
timestamp 1636968456
transform 1 0 58972 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_641
timestamp 1636968456
transform 1 0 60076 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_653
timestamp 1636968456
transform 1 0 61180 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_665
timestamp 1
transform 1 0 62284 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_671
timestamp 1
transform 1 0 62836 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_673
timestamp 1636968456
transform 1 0 63020 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_685
timestamp 1636968456
transform 1 0 64124 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_697
timestamp 1636968456
transform 1 0 65228 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_709
timestamp 1636968456
transform 1 0 66332 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_721
timestamp 1
transform 1 0 67436 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_727
timestamp 1
transform 1 0 67988 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_729
timestamp 1636968456
transform 1 0 68172 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_741
timestamp 1636968456
transform 1 0 69276 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_753
timestamp 1636968456
transform 1 0 70380 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_765
timestamp 1636968456
transform 1 0 71484 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_777
timestamp 1
transform 1 0 72588 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_783
timestamp 1
transform 1 0 73140 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_785
timestamp 1636968456
transform 1 0 73324 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_797
timestamp 1636968456
transform 1 0 74428 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_809
timestamp 1636968456
transform 1 0 75532 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_821
timestamp 1636968456
transform 1 0 76636 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_833
timestamp 1
transform 1 0 77740 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_839
timestamp 1
transform 1 0 78292 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_841
timestamp 1636968456
transform 1 0 78476 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_853
timestamp 1636968456
transform 1 0 79580 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_865
timestamp 1636968456
transform 1 0 80684 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_877
timestamp 1636968456
transform 1 0 81788 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_889
timestamp 1
transform 1 0 82892 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_895
timestamp 1
transform 1 0 83444 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_897
timestamp 1636968456
transform 1 0 83628 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_909
timestamp 1636968456
transform 1 0 84732 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_921
timestamp 1636968456
transform 1 0 85836 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_933
timestamp 1636968456
transform 1 0 86940 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_945
timestamp 1
transform 1 0 88044 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_951
timestamp 1
transform 1 0 88596 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_953
timestamp 1636968456
transform 1 0 88780 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_965
timestamp 1636968456
transform 1 0 89884 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_977
timestamp 1636968456
transform 1 0 90988 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_989
timestamp 1636968456
transform 1 0 92092 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_1001
timestamp 1
transform 1 0 93196 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_1007
timestamp 1
transform 1 0 93748 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_1009
timestamp 1636968456
transform 1 0 93932 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_1021
timestamp 1636968456
transform 1 0 95036 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_1033
timestamp 1636968456
transform 1 0 96140 0 -1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_113_1045
timestamp 1636968456
transform 1 0 97244 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_113_1057
timestamp 1
transform 1 0 98348 0 -1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_113_1063
timestamp 1
transform 1 0 98900 0 -1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_1065
timestamp 1636968456
transform 1 0 99084 0 -1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_113_1077
timestamp 1
transform 1 0 100188 0 -1 64192
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_114_3
timestamp 1636968456
transform 1 0 1380 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_15
timestamp 1636968456
transform 1 0 2484 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_114_27
timestamp 1
transform 1 0 3588 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_29
timestamp 1636968456
transform 1 0 3772 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_41
timestamp 1636968456
transform 1 0 4876 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_53
timestamp 1636968456
transform 1 0 5980 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_65
timestamp 1636968456
transform 1 0 7084 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_77
timestamp 1
transform 1 0 8188 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_83
timestamp 1
transform 1 0 8740 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_85
timestamp 1636968456
transform 1 0 8924 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_97
timestamp 1636968456
transform 1 0 10028 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_109
timestamp 1636968456
transform 1 0 11132 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_121
timestamp 1636968456
transform 1 0 12236 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_133
timestamp 1
transform 1 0 13340 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_139
timestamp 1
transform 1 0 13892 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_141
timestamp 1636968456
transform 1 0 14076 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_153
timestamp 1636968456
transform 1 0 15180 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_165
timestamp 1636968456
transform 1 0 16284 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_177
timestamp 1636968456
transform 1 0 17388 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_189
timestamp 1
transform 1 0 18492 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_195
timestamp 1
transform 1 0 19044 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_197
timestamp 1636968456
transform 1 0 19228 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_209
timestamp 1636968456
transform 1 0 20332 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_221
timestamp 1636968456
transform 1 0 21436 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_233
timestamp 1636968456
transform 1 0 22540 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_245
timestamp 1
transform 1 0 23644 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_251
timestamp 1
transform 1 0 24196 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_253
timestamp 1636968456
transform 1 0 24380 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_265
timestamp 1636968456
transform 1 0 25484 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_277
timestamp 1636968456
transform 1 0 26588 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_289
timestamp 1636968456
transform 1 0 27692 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_301
timestamp 1
transform 1 0 28796 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_307
timestamp 1
transform 1 0 29348 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_309
timestamp 1636968456
transform 1 0 29532 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_321
timestamp 1636968456
transform 1 0 30636 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_333
timestamp 1636968456
transform 1 0 31740 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_345
timestamp 1636968456
transform 1 0 32844 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_357
timestamp 1
transform 1 0 33948 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_363
timestamp 1
transform 1 0 34500 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_365
timestamp 1636968456
transform 1 0 34684 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_377
timestamp 1636968456
transform 1 0 35788 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_389
timestamp 1636968456
transform 1 0 36892 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_401
timestamp 1636968456
transform 1 0 37996 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_413
timestamp 1
transform 1 0 39100 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_419
timestamp 1
transform 1 0 39652 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_421
timestamp 1636968456
transform 1 0 39836 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_433
timestamp 1636968456
transform 1 0 40940 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_445
timestamp 1636968456
transform 1 0 42044 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_457
timestamp 1636968456
transform 1 0 43148 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_469
timestamp 1
transform 1 0 44252 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_475
timestamp 1
transform 1 0 44804 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_477
timestamp 1636968456
transform 1 0 44988 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_489
timestamp 1636968456
transform 1 0 46092 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_501
timestamp 1636968456
transform 1 0 47196 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_513
timestamp 1636968456
transform 1 0 48300 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_525
timestamp 1
transform 1 0 49404 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_531
timestamp 1
transform 1 0 49956 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_533
timestamp 1636968456
transform 1 0 50140 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_545
timestamp 1636968456
transform 1 0 51244 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_557
timestamp 1636968456
transform 1 0 52348 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_569
timestamp 1636968456
transform 1 0 53452 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_581
timestamp 1
transform 1 0 54556 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_587
timestamp 1
transform 1 0 55108 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_589
timestamp 1636968456
transform 1 0 55292 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_601
timestamp 1636968456
transform 1 0 56396 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_613
timestamp 1636968456
transform 1 0 57500 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_625
timestamp 1636968456
transform 1 0 58604 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_637
timestamp 1
transform 1 0 59708 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_643
timestamp 1
transform 1 0 60260 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_645
timestamp 1636968456
transform 1 0 60444 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_657
timestamp 1636968456
transform 1 0 61548 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_669
timestamp 1636968456
transform 1 0 62652 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_681
timestamp 1636968456
transform 1 0 63756 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_693
timestamp 1
transform 1 0 64860 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_699
timestamp 1
transform 1 0 65412 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_701
timestamp 1636968456
transform 1 0 65596 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_713
timestamp 1636968456
transform 1 0 66700 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_725
timestamp 1636968456
transform 1 0 67804 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_737
timestamp 1636968456
transform 1 0 68908 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_749
timestamp 1
transform 1 0 70012 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_755
timestamp 1
transform 1 0 70564 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_757
timestamp 1636968456
transform 1 0 70748 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_769
timestamp 1636968456
transform 1 0 71852 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_781
timestamp 1636968456
transform 1 0 72956 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_793
timestamp 1636968456
transform 1 0 74060 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_805
timestamp 1
transform 1 0 75164 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_811
timestamp 1
transform 1 0 75716 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_813
timestamp 1636968456
transform 1 0 75900 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_825
timestamp 1636968456
transform 1 0 77004 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_837
timestamp 1636968456
transform 1 0 78108 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_849
timestamp 1636968456
transform 1 0 79212 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_861
timestamp 1
transform 1 0 80316 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_867
timestamp 1
transform 1 0 80868 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_869
timestamp 1636968456
transform 1 0 81052 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_881
timestamp 1636968456
transform 1 0 82156 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_893
timestamp 1636968456
transform 1 0 83260 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_905
timestamp 1636968456
transform 1 0 84364 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_917
timestamp 1
transform 1 0 85468 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_923
timestamp 1
transform 1 0 86020 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_925
timestamp 1636968456
transform 1 0 86204 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_937
timestamp 1636968456
transform 1 0 87308 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_949
timestamp 1636968456
transform 1 0 88412 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_961
timestamp 1636968456
transform 1 0 89516 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_973
timestamp 1
transform 1 0 90620 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_979
timestamp 1
transform 1 0 91172 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_981
timestamp 1636968456
transform 1 0 91356 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_993
timestamp 1636968456
transform 1 0 92460 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_1005
timestamp 1636968456
transform 1 0 93564 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_1017
timestamp 1636968456
transform 1 0 94668 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_114_1029
timestamp 1
transform 1 0 95772 0 1 64192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_114_1035
timestamp 1
transform 1 0 96324 0 1 64192
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_1037
timestamp 1636968456
transform 1 0 96508 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_1049
timestamp 1636968456
transform 1 0 97612 0 1 64192
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_1061
timestamp 1636968456
transform 1 0 98716 0 1 64192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_114_1073
timestamp 1
transform 1 0 99820 0 1 64192
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_115_3
timestamp 1636968456
transform 1 0 1380 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_15
timestamp 1636968456
transform 1 0 2484 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_27
timestamp 1636968456
transform 1 0 3588 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_39
timestamp 1636968456
transform 1 0 4692 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_115_51
timestamp 1
transform 1 0 5796 0 -1 65280
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_115_55
timestamp 1
transform 1 0 6164 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_57
timestamp 1636968456
transform 1 0 6348 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_69
timestamp 1636968456
transform 1 0 7452 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_81
timestamp 1636968456
transform 1 0 8556 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_93
timestamp 1636968456
transform 1 0 9660 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_105
timestamp 1
transform 1 0 10764 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_111
timestamp 1
transform 1 0 11316 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_113
timestamp 1636968456
transform 1 0 11500 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_125
timestamp 1636968456
transform 1 0 12604 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_137
timestamp 1636968456
transform 1 0 13708 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_149
timestamp 1636968456
transform 1 0 14812 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_161
timestamp 1
transform 1 0 15916 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_167
timestamp 1
transform 1 0 16468 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_169
timestamp 1636968456
transform 1 0 16652 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_181
timestamp 1636968456
transform 1 0 17756 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_193
timestamp 1636968456
transform 1 0 18860 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_205
timestamp 1636968456
transform 1 0 19964 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_217
timestamp 1
transform 1 0 21068 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_223
timestamp 1
transform 1 0 21620 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_225
timestamp 1636968456
transform 1 0 21804 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_237
timestamp 1636968456
transform 1 0 22908 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_249
timestamp 1636968456
transform 1 0 24012 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_261
timestamp 1636968456
transform 1 0 25116 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_273
timestamp 1
transform 1 0 26220 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_279
timestamp 1
transform 1 0 26772 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_281
timestamp 1636968456
transform 1 0 26956 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_293
timestamp 1636968456
transform 1 0 28060 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_305
timestamp 1636968456
transform 1 0 29164 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_317
timestamp 1636968456
transform 1 0 30268 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_329
timestamp 1
transform 1 0 31372 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_335
timestamp 1
transform 1 0 31924 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_337
timestamp 1636968456
transform 1 0 32108 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_349
timestamp 1636968456
transform 1 0 33212 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_361
timestamp 1636968456
transform 1 0 34316 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_373
timestamp 1636968456
transform 1 0 35420 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_385
timestamp 1
transform 1 0 36524 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_391
timestamp 1
transform 1 0 37076 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_393
timestamp 1636968456
transform 1 0 37260 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_405
timestamp 1636968456
transform 1 0 38364 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_417
timestamp 1636968456
transform 1 0 39468 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_429
timestamp 1636968456
transform 1 0 40572 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_441
timestamp 1
transform 1 0 41676 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_447
timestamp 1
transform 1 0 42228 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_449
timestamp 1636968456
transform 1 0 42412 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_461
timestamp 1636968456
transform 1 0 43516 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_473
timestamp 1636968456
transform 1 0 44620 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_485
timestamp 1636968456
transform 1 0 45724 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_497
timestamp 1
transform 1 0 46828 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_503
timestamp 1
transform 1 0 47380 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_505
timestamp 1636968456
transform 1 0 47564 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_517
timestamp 1636968456
transform 1 0 48668 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_529
timestamp 1636968456
transform 1 0 49772 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_541
timestamp 1636968456
transform 1 0 50876 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_553
timestamp 1
transform 1 0 51980 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_559
timestamp 1
transform 1 0 52532 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_561
timestamp 1636968456
transform 1 0 52716 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_573
timestamp 1636968456
transform 1 0 53820 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_585
timestamp 1636968456
transform 1 0 54924 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_597
timestamp 1636968456
transform 1 0 56028 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_609
timestamp 1
transform 1 0 57132 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_615
timestamp 1
transform 1 0 57684 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_617
timestamp 1636968456
transform 1 0 57868 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_629
timestamp 1636968456
transform 1 0 58972 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_641
timestamp 1636968456
transform 1 0 60076 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_653
timestamp 1636968456
transform 1 0 61180 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_665
timestamp 1
transform 1 0 62284 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_671
timestamp 1
transform 1 0 62836 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_673
timestamp 1636968456
transform 1 0 63020 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_685
timestamp 1636968456
transform 1 0 64124 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_697
timestamp 1636968456
transform 1 0 65228 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_709
timestamp 1636968456
transform 1 0 66332 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_721
timestamp 1
transform 1 0 67436 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_727
timestamp 1
transform 1 0 67988 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_729
timestamp 1636968456
transform 1 0 68172 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_741
timestamp 1636968456
transform 1 0 69276 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_753
timestamp 1636968456
transform 1 0 70380 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_765
timestamp 1636968456
transform 1 0 71484 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_777
timestamp 1
transform 1 0 72588 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_783
timestamp 1
transform 1 0 73140 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_785
timestamp 1636968456
transform 1 0 73324 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_797
timestamp 1636968456
transform 1 0 74428 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_809
timestamp 1636968456
transform 1 0 75532 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_821
timestamp 1636968456
transform 1 0 76636 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_833
timestamp 1
transform 1 0 77740 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_839
timestamp 1
transform 1 0 78292 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_841
timestamp 1636968456
transform 1 0 78476 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_853
timestamp 1636968456
transform 1 0 79580 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_865
timestamp 1636968456
transform 1 0 80684 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_877
timestamp 1636968456
transform 1 0 81788 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_889
timestamp 1
transform 1 0 82892 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_895
timestamp 1
transform 1 0 83444 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_897
timestamp 1636968456
transform 1 0 83628 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_909
timestamp 1636968456
transform 1 0 84732 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_921
timestamp 1636968456
transform 1 0 85836 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_933
timestamp 1636968456
transform 1 0 86940 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_945
timestamp 1
transform 1 0 88044 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_951
timestamp 1
transform 1 0 88596 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_953
timestamp 1636968456
transform 1 0 88780 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_965
timestamp 1636968456
transform 1 0 89884 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_977
timestamp 1636968456
transform 1 0 90988 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_989
timestamp 1636968456
transform 1 0 92092 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_1001
timestamp 1
transform 1 0 93196 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_1007
timestamp 1
transform 1 0 93748 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_1009
timestamp 1636968456
transform 1 0 93932 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_1021
timestamp 1636968456
transform 1 0 95036 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_1033
timestamp 1636968456
transform 1 0 96140 0 -1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_115_1045
timestamp 1636968456
transform 1 0 97244 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_115_1057
timestamp 1
transform 1 0 98348 0 -1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_115_1063
timestamp 1
transform 1 0 98900 0 -1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_1065
timestamp 1636968456
transform 1 0 99084 0 -1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_115_1077
timestamp 1
transform 1 0 100188 0 -1 65280
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_116_3
timestamp 1636968456
transform 1 0 1380 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_15
timestamp 1636968456
transform 1 0 2484 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_116_27
timestamp 1
transform 1 0 3588 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_29
timestamp 1636968456
transform 1 0 3772 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_41
timestamp 1636968456
transform 1 0 4876 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_53
timestamp 1636968456
transform 1 0 5980 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_65
timestamp 1636968456
transform 1 0 7084 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_77
timestamp 1
transform 1 0 8188 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_83
timestamp 1
transform 1 0 8740 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_85
timestamp 1636968456
transform 1 0 8924 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_97
timestamp 1636968456
transform 1 0 10028 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_109
timestamp 1636968456
transform 1 0 11132 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_121
timestamp 1636968456
transform 1 0 12236 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_133
timestamp 1
transform 1 0 13340 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_139
timestamp 1
transform 1 0 13892 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_141
timestamp 1636968456
transform 1 0 14076 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_153
timestamp 1636968456
transform 1 0 15180 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_165
timestamp 1636968456
transform 1 0 16284 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_177
timestamp 1636968456
transform 1 0 17388 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_189
timestamp 1
transform 1 0 18492 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_195
timestamp 1
transform 1 0 19044 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_197
timestamp 1636968456
transform 1 0 19228 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_209
timestamp 1636968456
transform 1 0 20332 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_221
timestamp 1636968456
transform 1 0 21436 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_233
timestamp 1636968456
transform 1 0 22540 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_245
timestamp 1
transform 1 0 23644 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_251
timestamp 1
transform 1 0 24196 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_253
timestamp 1636968456
transform 1 0 24380 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_265
timestamp 1636968456
transform 1 0 25484 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_277
timestamp 1636968456
transform 1 0 26588 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_289
timestamp 1636968456
transform 1 0 27692 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_301
timestamp 1
transform 1 0 28796 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_307
timestamp 1
transform 1 0 29348 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_309
timestamp 1636968456
transform 1 0 29532 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_321
timestamp 1636968456
transform 1 0 30636 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_333
timestamp 1636968456
transform 1 0 31740 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_345
timestamp 1636968456
transform 1 0 32844 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_357
timestamp 1
transform 1 0 33948 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_363
timestamp 1
transform 1 0 34500 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_365
timestamp 1636968456
transform 1 0 34684 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_377
timestamp 1636968456
transform 1 0 35788 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_389
timestamp 1636968456
transform 1 0 36892 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_401
timestamp 1636968456
transform 1 0 37996 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_413
timestamp 1
transform 1 0 39100 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_419
timestamp 1
transform 1 0 39652 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_421
timestamp 1636968456
transform 1 0 39836 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_433
timestamp 1636968456
transform 1 0 40940 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_445
timestamp 1636968456
transform 1 0 42044 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_457
timestamp 1636968456
transform 1 0 43148 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_469
timestamp 1
transform 1 0 44252 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_475
timestamp 1
transform 1 0 44804 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_477
timestamp 1636968456
transform 1 0 44988 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_489
timestamp 1636968456
transform 1 0 46092 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_501
timestamp 1636968456
transform 1 0 47196 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_513
timestamp 1636968456
transform 1 0 48300 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_525
timestamp 1
transform 1 0 49404 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_531
timestamp 1
transform 1 0 49956 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_533
timestamp 1636968456
transform 1 0 50140 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_545
timestamp 1636968456
transform 1 0 51244 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_557
timestamp 1636968456
transform 1 0 52348 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_569
timestamp 1636968456
transform 1 0 53452 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_581
timestamp 1
transform 1 0 54556 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_587
timestamp 1
transform 1 0 55108 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_589
timestamp 1636968456
transform 1 0 55292 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_601
timestamp 1636968456
transform 1 0 56396 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_613
timestamp 1636968456
transform 1 0 57500 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_625
timestamp 1636968456
transform 1 0 58604 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_637
timestamp 1
transform 1 0 59708 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_643
timestamp 1
transform 1 0 60260 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_645
timestamp 1636968456
transform 1 0 60444 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_657
timestamp 1636968456
transform 1 0 61548 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_669
timestamp 1636968456
transform 1 0 62652 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_681
timestamp 1636968456
transform 1 0 63756 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_693
timestamp 1
transform 1 0 64860 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_699
timestamp 1
transform 1 0 65412 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_701
timestamp 1636968456
transform 1 0 65596 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_713
timestamp 1636968456
transform 1 0 66700 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_725
timestamp 1636968456
transform 1 0 67804 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_737
timestamp 1636968456
transform 1 0 68908 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_749
timestamp 1
transform 1 0 70012 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_755
timestamp 1
transform 1 0 70564 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_757
timestamp 1636968456
transform 1 0 70748 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_769
timestamp 1636968456
transform 1 0 71852 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_781
timestamp 1636968456
transform 1 0 72956 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_793
timestamp 1636968456
transform 1 0 74060 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_805
timestamp 1
transform 1 0 75164 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_811
timestamp 1
transform 1 0 75716 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_813
timestamp 1636968456
transform 1 0 75900 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_825
timestamp 1636968456
transform 1 0 77004 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_837
timestamp 1636968456
transform 1 0 78108 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_849
timestamp 1636968456
transform 1 0 79212 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_861
timestamp 1
transform 1 0 80316 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_867
timestamp 1
transform 1 0 80868 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_869
timestamp 1636968456
transform 1 0 81052 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_881
timestamp 1636968456
transform 1 0 82156 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_893
timestamp 1636968456
transform 1 0 83260 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_905
timestamp 1636968456
transform 1 0 84364 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_917
timestamp 1
transform 1 0 85468 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_923
timestamp 1
transform 1 0 86020 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_925
timestamp 1636968456
transform 1 0 86204 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_937
timestamp 1636968456
transform 1 0 87308 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_949
timestamp 1636968456
transform 1 0 88412 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_961
timestamp 1636968456
transform 1 0 89516 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_973
timestamp 1
transform 1 0 90620 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_979
timestamp 1
transform 1 0 91172 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_981
timestamp 1636968456
transform 1 0 91356 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_993
timestamp 1636968456
transform 1 0 92460 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_1005
timestamp 1636968456
transform 1 0 93564 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_1017
timestamp 1636968456
transform 1 0 94668 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_116_1029
timestamp 1
transform 1 0 95772 0 1 65280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_116_1035
timestamp 1
transform 1 0 96324 0 1 65280
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_1037
timestamp 1636968456
transform 1 0 96508 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_1049
timestamp 1636968456
transform 1 0 97612 0 1 65280
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_1061
timestamp 1636968456
transform 1 0 98716 0 1 65280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_116_1073
timestamp 1
transform 1 0 99820 0 1 65280
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_117_3
timestamp 1636968456
transform 1 0 1380 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_15
timestamp 1636968456
transform 1 0 2484 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_27
timestamp 1636968456
transform 1 0 3588 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_39
timestamp 1636968456
transform 1 0 4692 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_117_51
timestamp 1
transform 1 0 5796 0 -1 66368
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_117_55
timestamp 1
transform 1 0 6164 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_57
timestamp 1636968456
transform 1 0 6348 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_69
timestamp 1636968456
transform 1 0 7452 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_81
timestamp 1636968456
transform 1 0 8556 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_93
timestamp 1636968456
transform 1 0 9660 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_105
timestamp 1
transform 1 0 10764 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_111
timestamp 1
transform 1 0 11316 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_113
timestamp 1636968456
transform 1 0 11500 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_125
timestamp 1636968456
transform 1 0 12604 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_137
timestamp 1636968456
transform 1 0 13708 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_149
timestamp 1636968456
transform 1 0 14812 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_161
timestamp 1
transform 1 0 15916 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_167
timestamp 1
transform 1 0 16468 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_169
timestamp 1636968456
transform 1 0 16652 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_181
timestamp 1636968456
transform 1 0 17756 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_193
timestamp 1636968456
transform 1 0 18860 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_205
timestamp 1636968456
transform 1 0 19964 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_217
timestamp 1
transform 1 0 21068 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_223
timestamp 1
transform 1 0 21620 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_225
timestamp 1636968456
transform 1 0 21804 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_237
timestamp 1636968456
transform 1 0 22908 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_249
timestamp 1636968456
transform 1 0 24012 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_261
timestamp 1636968456
transform 1 0 25116 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_273
timestamp 1
transform 1 0 26220 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_279
timestamp 1
transform 1 0 26772 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_281
timestamp 1636968456
transform 1 0 26956 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_293
timestamp 1636968456
transform 1 0 28060 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_305
timestamp 1636968456
transform 1 0 29164 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_317
timestamp 1636968456
transform 1 0 30268 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_329
timestamp 1
transform 1 0 31372 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_335
timestamp 1
transform 1 0 31924 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_337
timestamp 1636968456
transform 1 0 32108 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_349
timestamp 1636968456
transform 1 0 33212 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_361
timestamp 1636968456
transform 1 0 34316 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_373
timestamp 1636968456
transform 1 0 35420 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_385
timestamp 1
transform 1 0 36524 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_391
timestamp 1
transform 1 0 37076 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_393
timestamp 1636968456
transform 1 0 37260 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_405
timestamp 1636968456
transform 1 0 38364 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_417
timestamp 1636968456
transform 1 0 39468 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_429
timestamp 1636968456
transform 1 0 40572 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_441
timestamp 1
transform 1 0 41676 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_447
timestamp 1
transform 1 0 42228 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_449
timestamp 1636968456
transform 1 0 42412 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_461
timestamp 1636968456
transform 1 0 43516 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_473
timestamp 1636968456
transform 1 0 44620 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_485
timestamp 1636968456
transform 1 0 45724 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_497
timestamp 1
transform 1 0 46828 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_503
timestamp 1
transform 1 0 47380 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_505
timestamp 1636968456
transform 1 0 47564 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_517
timestamp 1636968456
transform 1 0 48668 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_529
timestamp 1636968456
transform 1 0 49772 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_541
timestamp 1636968456
transform 1 0 50876 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_553
timestamp 1
transform 1 0 51980 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_559
timestamp 1
transform 1 0 52532 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_561
timestamp 1636968456
transform 1 0 52716 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_573
timestamp 1636968456
transform 1 0 53820 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_585
timestamp 1636968456
transform 1 0 54924 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_597
timestamp 1636968456
transform 1 0 56028 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_609
timestamp 1
transform 1 0 57132 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_615
timestamp 1
transform 1 0 57684 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_617
timestamp 1636968456
transform 1 0 57868 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_629
timestamp 1636968456
transform 1 0 58972 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_641
timestamp 1636968456
transform 1 0 60076 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_653
timestamp 1636968456
transform 1 0 61180 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_665
timestamp 1
transform 1 0 62284 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_671
timestamp 1
transform 1 0 62836 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_673
timestamp 1636968456
transform 1 0 63020 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_685
timestamp 1636968456
transform 1 0 64124 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_697
timestamp 1636968456
transform 1 0 65228 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_709
timestamp 1636968456
transform 1 0 66332 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_721
timestamp 1
transform 1 0 67436 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_727
timestamp 1
transform 1 0 67988 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_729
timestamp 1636968456
transform 1 0 68172 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_741
timestamp 1636968456
transform 1 0 69276 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_753
timestamp 1636968456
transform 1 0 70380 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_765
timestamp 1636968456
transform 1 0 71484 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_777
timestamp 1
transform 1 0 72588 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_783
timestamp 1
transform 1 0 73140 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_785
timestamp 1636968456
transform 1 0 73324 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_797
timestamp 1636968456
transform 1 0 74428 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_809
timestamp 1636968456
transform 1 0 75532 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_821
timestamp 1636968456
transform 1 0 76636 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_833
timestamp 1
transform 1 0 77740 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_839
timestamp 1
transform 1 0 78292 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_841
timestamp 1636968456
transform 1 0 78476 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_853
timestamp 1636968456
transform 1 0 79580 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_865
timestamp 1636968456
transform 1 0 80684 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_877
timestamp 1636968456
transform 1 0 81788 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_889
timestamp 1
transform 1 0 82892 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_895
timestamp 1
transform 1 0 83444 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_897
timestamp 1636968456
transform 1 0 83628 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_909
timestamp 1636968456
transform 1 0 84732 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_921
timestamp 1636968456
transform 1 0 85836 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_933
timestamp 1636968456
transform 1 0 86940 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_945
timestamp 1
transform 1 0 88044 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_951
timestamp 1
transform 1 0 88596 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_953
timestamp 1636968456
transform 1 0 88780 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_965
timestamp 1636968456
transform 1 0 89884 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_977
timestamp 1636968456
transform 1 0 90988 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_989
timestamp 1636968456
transform 1 0 92092 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_1001
timestamp 1
transform 1 0 93196 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_1007
timestamp 1
transform 1 0 93748 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_1009
timestamp 1636968456
transform 1 0 93932 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_1021
timestamp 1636968456
transform 1 0 95036 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_1033
timestamp 1636968456
transform 1 0 96140 0 -1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_117_1045
timestamp 1636968456
transform 1 0 97244 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_117_1057
timestamp 1
transform 1 0 98348 0 -1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_117_1063
timestamp 1
transform 1 0 98900 0 -1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_1065
timestamp 1636968456
transform 1 0 99084 0 -1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_117_1077
timestamp 1
transform 1 0 100188 0 -1 66368
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_118_3
timestamp 1636968456
transform 1 0 1380 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_15
timestamp 1636968456
transform 1 0 2484 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_118_27
timestamp 1
transform 1 0 3588 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_29
timestamp 1636968456
transform 1 0 3772 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_41
timestamp 1636968456
transform 1 0 4876 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_53
timestamp 1636968456
transform 1 0 5980 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_65
timestamp 1636968456
transform 1 0 7084 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_77
timestamp 1
transform 1 0 8188 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_83
timestamp 1
transform 1 0 8740 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_85
timestamp 1636968456
transform 1 0 8924 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_97
timestamp 1636968456
transform 1 0 10028 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_109
timestamp 1636968456
transform 1 0 11132 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_121
timestamp 1636968456
transform 1 0 12236 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_133
timestamp 1
transform 1 0 13340 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_139
timestamp 1
transform 1 0 13892 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_141
timestamp 1636968456
transform 1 0 14076 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_153
timestamp 1636968456
transform 1 0 15180 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_165
timestamp 1636968456
transform 1 0 16284 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_177
timestamp 1636968456
transform 1 0 17388 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_189
timestamp 1
transform 1 0 18492 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_195
timestamp 1
transform 1 0 19044 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_197
timestamp 1636968456
transform 1 0 19228 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_209
timestamp 1636968456
transform 1 0 20332 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_221
timestamp 1636968456
transform 1 0 21436 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_233
timestamp 1636968456
transform 1 0 22540 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_245
timestamp 1
transform 1 0 23644 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_251
timestamp 1
transform 1 0 24196 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_253
timestamp 1636968456
transform 1 0 24380 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_265
timestamp 1636968456
transform 1 0 25484 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_277
timestamp 1636968456
transform 1 0 26588 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_289
timestamp 1636968456
transform 1 0 27692 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_301
timestamp 1
transform 1 0 28796 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_307
timestamp 1
transform 1 0 29348 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_309
timestamp 1636968456
transform 1 0 29532 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_321
timestamp 1636968456
transform 1 0 30636 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_333
timestamp 1636968456
transform 1 0 31740 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_345
timestamp 1636968456
transform 1 0 32844 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_357
timestamp 1
transform 1 0 33948 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_363
timestamp 1
transform 1 0 34500 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_365
timestamp 1636968456
transform 1 0 34684 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_377
timestamp 1636968456
transform 1 0 35788 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_389
timestamp 1636968456
transform 1 0 36892 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_401
timestamp 1636968456
transform 1 0 37996 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_413
timestamp 1
transform 1 0 39100 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_419
timestamp 1
transform 1 0 39652 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_421
timestamp 1636968456
transform 1 0 39836 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_433
timestamp 1636968456
transform 1 0 40940 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_445
timestamp 1636968456
transform 1 0 42044 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_457
timestamp 1636968456
transform 1 0 43148 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_469
timestamp 1
transform 1 0 44252 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_475
timestamp 1
transform 1 0 44804 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_477
timestamp 1636968456
transform 1 0 44988 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_489
timestamp 1636968456
transform 1 0 46092 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_501
timestamp 1636968456
transform 1 0 47196 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_513
timestamp 1636968456
transform 1 0 48300 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_525
timestamp 1
transform 1 0 49404 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_531
timestamp 1
transform 1 0 49956 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_533
timestamp 1636968456
transform 1 0 50140 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_545
timestamp 1636968456
transform 1 0 51244 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_557
timestamp 1636968456
transform 1 0 52348 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_569
timestamp 1636968456
transform 1 0 53452 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_581
timestamp 1
transform 1 0 54556 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_587
timestamp 1
transform 1 0 55108 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_589
timestamp 1636968456
transform 1 0 55292 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_601
timestamp 1636968456
transform 1 0 56396 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_613
timestamp 1636968456
transform 1 0 57500 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_625
timestamp 1636968456
transform 1 0 58604 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_637
timestamp 1
transform 1 0 59708 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_643
timestamp 1
transform 1 0 60260 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_645
timestamp 1636968456
transform 1 0 60444 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_657
timestamp 1636968456
transform 1 0 61548 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_669
timestamp 1636968456
transform 1 0 62652 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_681
timestamp 1636968456
transform 1 0 63756 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_693
timestamp 1
transform 1 0 64860 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_699
timestamp 1
transform 1 0 65412 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_701
timestamp 1636968456
transform 1 0 65596 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_713
timestamp 1636968456
transform 1 0 66700 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_725
timestamp 1636968456
transform 1 0 67804 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_737
timestamp 1636968456
transform 1 0 68908 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_749
timestamp 1
transform 1 0 70012 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_755
timestamp 1
transform 1 0 70564 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_757
timestamp 1636968456
transform 1 0 70748 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_769
timestamp 1636968456
transform 1 0 71852 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_781
timestamp 1636968456
transform 1 0 72956 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_793
timestamp 1636968456
transform 1 0 74060 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_805
timestamp 1
transform 1 0 75164 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_811
timestamp 1
transform 1 0 75716 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_813
timestamp 1636968456
transform 1 0 75900 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_825
timestamp 1636968456
transform 1 0 77004 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_837
timestamp 1636968456
transform 1 0 78108 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_849
timestamp 1636968456
transform 1 0 79212 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_861
timestamp 1
transform 1 0 80316 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_867
timestamp 1
transform 1 0 80868 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_869
timestamp 1636968456
transform 1 0 81052 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_881
timestamp 1636968456
transform 1 0 82156 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_893
timestamp 1636968456
transform 1 0 83260 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_905
timestamp 1636968456
transform 1 0 84364 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_917
timestamp 1
transform 1 0 85468 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_923
timestamp 1
transform 1 0 86020 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_925
timestamp 1636968456
transform 1 0 86204 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_937
timestamp 1636968456
transform 1 0 87308 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_949
timestamp 1636968456
transform 1 0 88412 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_961
timestamp 1636968456
transform 1 0 89516 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_973
timestamp 1
transform 1 0 90620 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_979
timestamp 1
transform 1 0 91172 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_981
timestamp 1636968456
transform 1 0 91356 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_993
timestamp 1636968456
transform 1 0 92460 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_1005
timestamp 1636968456
transform 1 0 93564 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_1017
timestamp 1636968456
transform 1 0 94668 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_118_1029
timestamp 1
transform 1 0 95772 0 1 66368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_118_1035
timestamp 1
transform 1 0 96324 0 1 66368
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_1037
timestamp 1636968456
transform 1 0 96508 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_1049
timestamp 1636968456
transform 1 0 97612 0 1 66368
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_1061
timestamp 1636968456
transform 1 0 98716 0 1 66368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_118_1073
timestamp 1
transform 1 0 99820 0 1 66368
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_119_3
timestamp 1636968456
transform 1 0 1380 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_15
timestamp 1636968456
transform 1 0 2484 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_27
timestamp 1636968456
transform 1 0 3588 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_39
timestamp 1636968456
transform 1 0 4692 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_119_51
timestamp 1
transform 1 0 5796 0 -1 67456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_119_55
timestamp 1
transform 1 0 6164 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_57
timestamp 1636968456
transform 1 0 6348 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_69
timestamp 1636968456
transform 1 0 7452 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_81
timestamp 1636968456
transform 1 0 8556 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_93
timestamp 1636968456
transform 1 0 9660 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_105
timestamp 1
transform 1 0 10764 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_111
timestamp 1
transform 1 0 11316 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_113
timestamp 1636968456
transform 1 0 11500 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_125
timestamp 1636968456
transform 1 0 12604 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_137
timestamp 1636968456
transform 1 0 13708 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_149
timestamp 1636968456
transform 1 0 14812 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_161
timestamp 1
transform 1 0 15916 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_167
timestamp 1
transform 1 0 16468 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_169
timestamp 1636968456
transform 1 0 16652 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_181
timestamp 1636968456
transform 1 0 17756 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_193
timestamp 1636968456
transform 1 0 18860 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_205
timestamp 1636968456
transform 1 0 19964 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_217
timestamp 1
transform 1 0 21068 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_223
timestamp 1
transform 1 0 21620 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_225
timestamp 1636968456
transform 1 0 21804 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_237
timestamp 1636968456
transform 1 0 22908 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_249
timestamp 1636968456
transform 1 0 24012 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_261
timestamp 1636968456
transform 1 0 25116 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_273
timestamp 1
transform 1 0 26220 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_279
timestamp 1
transform 1 0 26772 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_281
timestamp 1636968456
transform 1 0 26956 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_293
timestamp 1636968456
transform 1 0 28060 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_305
timestamp 1636968456
transform 1 0 29164 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_317
timestamp 1636968456
transform 1 0 30268 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_329
timestamp 1
transform 1 0 31372 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_335
timestamp 1
transform 1 0 31924 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_337
timestamp 1636968456
transform 1 0 32108 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_349
timestamp 1636968456
transform 1 0 33212 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_361
timestamp 1636968456
transform 1 0 34316 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_373
timestamp 1636968456
transform 1 0 35420 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_385
timestamp 1
transform 1 0 36524 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_391
timestamp 1
transform 1 0 37076 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_393
timestamp 1636968456
transform 1 0 37260 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_405
timestamp 1636968456
transform 1 0 38364 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_417
timestamp 1636968456
transform 1 0 39468 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_429
timestamp 1636968456
transform 1 0 40572 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_441
timestamp 1
transform 1 0 41676 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_447
timestamp 1
transform 1 0 42228 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_449
timestamp 1636968456
transform 1 0 42412 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_461
timestamp 1636968456
transform 1 0 43516 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_473
timestamp 1636968456
transform 1 0 44620 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_485
timestamp 1636968456
transform 1 0 45724 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_497
timestamp 1
transform 1 0 46828 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_503
timestamp 1
transform 1 0 47380 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_505
timestamp 1636968456
transform 1 0 47564 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_517
timestamp 1636968456
transform 1 0 48668 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_529
timestamp 1636968456
transform 1 0 49772 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_541
timestamp 1636968456
transform 1 0 50876 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_553
timestamp 1
transform 1 0 51980 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_559
timestamp 1
transform 1 0 52532 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_561
timestamp 1636968456
transform 1 0 52716 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_573
timestamp 1636968456
transform 1 0 53820 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_585
timestamp 1636968456
transform 1 0 54924 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_597
timestamp 1636968456
transform 1 0 56028 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_609
timestamp 1
transform 1 0 57132 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_615
timestamp 1
transform 1 0 57684 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_617
timestamp 1636968456
transform 1 0 57868 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_629
timestamp 1636968456
transform 1 0 58972 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_641
timestamp 1636968456
transform 1 0 60076 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_653
timestamp 1636968456
transform 1 0 61180 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_665
timestamp 1
transform 1 0 62284 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_671
timestamp 1
transform 1 0 62836 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_673
timestamp 1636968456
transform 1 0 63020 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_685
timestamp 1636968456
transform 1 0 64124 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_697
timestamp 1636968456
transform 1 0 65228 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_709
timestamp 1636968456
transform 1 0 66332 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_721
timestamp 1
transform 1 0 67436 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_727
timestamp 1
transform 1 0 67988 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_729
timestamp 1636968456
transform 1 0 68172 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_741
timestamp 1636968456
transform 1 0 69276 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_753
timestamp 1636968456
transform 1 0 70380 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_765
timestamp 1636968456
transform 1 0 71484 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_777
timestamp 1
transform 1 0 72588 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_783
timestamp 1
transform 1 0 73140 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_785
timestamp 1636968456
transform 1 0 73324 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_797
timestamp 1636968456
transform 1 0 74428 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_809
timestamp 1636968456
transform 1 0 75532 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_821
timestamp 1636968456
transform 1 0 76636 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_833
timestamp 1
transform 1 0 77740 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_839
timestamp 1
transform 1 0 78292 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_841
timestamp 1636968456
transform 1 0 78476 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_853
timestamp 1636968456
transform 1 0 79580 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_865
timestamp 1636968456
transform 1 0 80684 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_877
timestamp 1636968456
transform 1 0 81788 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_889
timestamp 1
transform 1 0 82892 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_895
timestamp 1
transform 1 0 83444 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_897
timestamp 1636968456
transform 1 0 83628 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_909
timestamp 1636968456
transform 1 0 84732 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_921
timestamp 1636968456
transform 1 0 85836 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_933
timestamp 1636968456
transform 1 0 86940 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_945
timestamp 1
transform 1 0 88044 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_951
timestamp 1
transform 1 0 88596 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_953
timestamp 1636968456
transform 1 0 88780 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_965
timestamp 1636968456
transform 1 0 89884 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_977
timestamp 1636968456
transform 1 0 90988 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_989
timestamp 1636968456
transform 1 0 92092 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_1001
timestamp 1
transform 1 0 93196 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_1007
timestamp 1
transform 1 0 93748 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_1009
timestamp 1636968456
transform 1 0 93932 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_1021
timestamp 1636968456
transform 1 0 95036 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_1033
timestamp 1636968456
transform 1 0 96140 0 -1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_119_1045
timestamp 1636968456
transform 1 0 97244 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_1057
timestamp 1
transform 1 0 98348 0 -1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_119_1063
timestamp 1
transform 1 0 98900 0 -1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_119_1065
timestamp 1636968456
transform 1 0 99084 0 -1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_119_1077
timestamp 1
transform 1 0 100188 0 -1 67456
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_120_3
timestamp 1636968456
transform 1 0 1380 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_15
timestamp 1636968456
transform 1 0 2484 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_120_27
timestamp 1
transform 1 0 3588 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_29
timestamp 1636968456
transform 1 0 3772 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_41
timestamp 1636968456
transform 1 0 4876 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_53
timestamp 1636968456
transform 1 0 5980 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_65
timestamp 1636968456
transform 1 0 7084 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_77
timestamp 1
transform 1 0 8188 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_83
timestamp 1
transform 1 0 8740 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_85
timestamp 1636968456
transform 1 0 8924 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_97
timestamp 1636968456
transform 1 0 10028 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_109
timestamp 1636968456
transform 1 0 11132 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_121
timestamp 1636968456
transform 1 0 12236 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_133
timestamp 1
transform 1 0 13340 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_139
timestamp 1
transform 1 0 13892 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_141
timestamp 1636968456
transform 1 0 14076 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_153
timestamp 1636968456
transform 1 0 15180 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_165
timestamp 1636968456
transform 1 0 16284 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_177
timestamp 1636968456
transform 1 0 17388 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_189
timestamp 1
transform 1 0 18492 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_195
timestamp 1
transform 1 0 19044 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_197
timestamp 1636968456
transform 1 0 19228 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_209
timestamp 1636968456
transform 1 0 20332 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_221
timestamp 1636968456
transform 1 0 21436 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_233
timestamp 1636968456
transform 1 0 22540 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_245
timestamp 1
transform 1 0 23644 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_251
timestamp 1
transform 1 0 24196 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_253
timestamp 1636968456
transform 1 0 24380 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_265
timestamp 1636968456
transform 1 0 25484 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_277
timestamp 1636968456
transform 1 0 26588 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_289
timestamp 1636968456
transform 1 0 27692 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_301
timestamp 1
transform 1 0 28796 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_307
timestamp 1
transform 1 0 29348 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_309
timestamp 1636968456
transform 1 0 29532 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_321
timestamp 1636968456
transform 1 0 30636 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_333
timestamp 1636968456
transform 1 0 31740 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_345
timestamp 1636968456
transform 1 0 32844 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_357
timestamp 1
transform 1 0 33948 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_363
timestamp 1
transform 1 0 34500 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_365
timestamp 1636968456
transform 1 0 34684 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_377
timestamp 1636968456
transform 1 0 35788 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_389
timestamp 1636968456
transform 1 0 36892 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_401
timestamp 1636968456
transform 1 0 37996 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_413
timestamp 1
transform 1 0 39100 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_419
timestamp 1
transform 1 0 39652 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_421
timestamp 1636968456
transform 1 0 39836 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_433
timestamp 1636968456
transform 1 0 40940 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_445
timestamp 1636968456
transform 1 0 42044 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_457
timestamp 1636968456
transform 1 0 43148 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_469
timestamp 1
transform 1 0 44252 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_475
timestamp 1
transform 1 0 44804 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_477
timestamp 1636968456
transform 1 0 44988 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_489
timestamp 1636968456
transform 1 0 46092 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_501
timestamp 1636968456
transform 1 0 47196 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_513
timestamp 1636968456
transform 1 0 48300 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_525
timestamp 1
transform 1 0 49404 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_531
timestamp 1
transform 1 0 49956 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_533
timestamp 1636968456
transform 1 0 50140 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_545
timestamp 1636968456
transform 1 0 51244 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_557
timestamp 1636968456
transform 1 0 52348 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_569
timestamp 1636968456
transform 1 0 53452 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_581
timestamp 1
transform 1 0 54556 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_587
timestamp 1
transform 1 0 55108 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_589
timestamp 1636968456
transform 1 0 55292 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_601
timestamp 1636968456
transform 1 0 56396 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_613
timestamp 1636968456
transform 1 0 57500 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_625
timestamp 1636968456
transform 1 0 58604 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_637
timestamp 1
transform 1 0 59708 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_643
timestamp 1
transform 1 0 60260 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_645
timestamp 1636968456
transform 1 0 60444 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_657
timestamp 1636968456
transform 1 0 61548 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_669
timestamp 1636968456
transform 1 0 62652 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_681
timestamp 1636968456
transform 1 0 63756 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_693
timestamp 1
transform 1 0 64860 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_699
timestamp 1
transform 1 0 65412 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_701
timestamp 1636968456
transform 1 0 65596 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_713
timestamp 1636968456
transform 1 0 66700 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_725
timestamp 1636968456
transform 1 0 67804 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_737
timestamp 1636968456
transform 1 0 68908 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_749
timestamp 1
transform 1 0 70012 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_755
timestamp 1
transform 1 0 70564 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_757
timestamp 1636968456
transform 1 0 70748 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_769
timestamp 1636968456
transform 1 0 71852 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_781
timestamp 1636968456
transform 1 0 72956 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_793
timestamp 1636968456
transform 1 0 74060 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_805
timestamp 1
transform 1 0 75164 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_811
timestamp 1
transform 1 0 75716 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_813
timestamp 1636968456
transform 1 0 75900 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_825
timestamp 1636968456
transform 1 0 77004 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_837
timestamp 1636968456
transform 1 0 78108 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_849
timestamp 1636968456
transform 1 0 79212 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_861
timestamp 1
transform 1 0 80316 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_867
timestamp 1
transform 1 0 80868 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_869
timestamp 1636968456
transform 1 0 81052 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_881
timestamp 1636968456
transform 1 0 82156 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_893
timestamp 1636968456
transform 1 0 83260 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_905
timestamp 1636968456
transform 1 0 84364 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_917
timestamp 1
transform 1 0 85468 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_923
timestamp 1
transform 1 0 86020 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_925
timestamp 1636968456
transform 1 0 86204 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_937
timestamp 1636968456
transform 1 0 87308 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_949
timestamp 1636968456
transform 1 0 88412 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_961
timestamp 1636968456
transform 1 0 89516 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_973
timestamp 1
transform 1 0 90620 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_979
timestamp 1
transform 1 0 91172 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_981
timestamp 1636968456
transform 1 0 91356 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_993
timestamp 1636968456
transform 1 0 92460 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_1005
timestamp 1636968456
transform 1 0 93564 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_1017
timestamp 1636968456
transform 1 0 94668 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_120_1029
timestamp 1
transform 1 0 95772 0 1 67456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_120_1035
timestamp 1
transform 1 0 96324 0 1 67456
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_1037
timestamp 1636968456
transform 1 0 96508 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_1049
timestamp 1636968456
transform 1 0 97612 0 1 67456
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_120_1061
timestamp 1636968456
transform 1 0 98716 0 1 67456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_120_1073
timestamp 1
transform 1 0 99820 0 1 67456
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_121_3
timestamp 1636968456
transform 1 0 1380 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_15
timestamp 1636968456
transform 1 0 2484 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_27
timestamp 1636968456
transform 1 0 3588 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_39
timestamp 1636968456
transform 1 0 4692 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_121_51
timestamp 1
transform 1 0 5796 0 -1 68544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_121_55
timestamp 1
transform 1 0 6164 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_57
timestamp 1636968456
transform 1 0 6348 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_69
timestamp 1636968456
transform 1 0 7452 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_81
timestamp 1636968456
transform 1 0 8556 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_93
timestamp 1636968456
transform 1 0 9660 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_105
timestamp 1
transform 1 0 10764 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_111
timestamp 1
transform 1 0 11316 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_113
timestamp 1636968456
transform 1 0 11500 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_125
timestamp 1636968456
transform 1 0 12604 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_137
timestamp 1636968456
transform 1 0 13708 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_149
timestamp 1636968456
transform 1 0 14812 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_161
timestamp 1
transform 1 0 15916 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_167
timestamp 1
transform 1 0 16468 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_169
timestamp 1636968456
transform 1 0 16652 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_181
timestamp 1636968456
transform 1 0 17756 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_193
timestamp 1636968456
transform 1 0 18860 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_205
timestamp 1636968456
transform 1 0 19964 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_217
timestamp 1
transform 1 0 21068 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_223
timestamp 1
transform 1 0 21620 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_225
timestamp 1636968456
transform 1 0 21804 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_237
timestamp 1636968456
transform 1 0 22908 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_249
timestamp 1636968456
transform 1 0 24012 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_261
timestamp 1636968456
transform 1 0 25116 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_273
timestamp 1
transform 1 0 26220 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_279
timestamp 1
transform 1 0 26772 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_281
timestamp 1636968456
transform 1 0 26956 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_293
timestamp 1636968456
transform 1 0 28060 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_305
timestamp 1636968456
transform 1 0 29164 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_317
timestamp 1636968456
transform 1 0 30268 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_329
timestamp 1
transform 1 0 31372 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_335
timestamp 1
transform 1 0 31924 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_337
timestamp 1636968456
transform 1 0 32108 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_349
timestamp 1636968456
transform 1 0 33212 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_361
timestamp 1636968456
transform 1 0 34316 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_373
timestamp 1636968456
transform 1 0 35420 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_385
timestamp 1
transform 1 0 36524 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_391
timestamp 1
transform 1 0 37076 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_393
timestamp 1636968456
transform 1 0 37260 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_405
timestamp 1636968456
transform 1 0 38364 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_417
timestamp 1636968456
transform 1 0 39468 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_429
timestamp 1636968456
transform 1 0 40572 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_441
timestamp 1
transform 1 0 41676 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_447
timestamp 1
transform 1 0 42228 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_449
timestamp 1636968456
transform 1 0 42412 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_461
timestamp 1636968456
transform 1 0 43516 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_473
timestamp 1636968456
transform 1 0 44620 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_485
timestamp 1636968456
transform 1 0 45724 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_497
timestamp 1
transform 1 0 46828 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_503
timestamp 1
transform 1 0 47380 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_505
timestamp 1636968456
transform 1 0 47564 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_517
timestamp 1636968456
transform 1 0 48668 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_529
timestamp 1636968456
transform 1 0 49772 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_541
timestamp 1636968456
transform 1 0 50876 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_553
timestamp 1
transform 1 0 51980 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_559
timestamp 1
transform 1 0 52532 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_561
timestamp 1636968456
transform 1 0 52716 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_573
timestamp 1636968456
transform 1 0 53820 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_585
timestamp 1636968456
transform 1 0 54924 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_597
timestamp 1636968456
transform 1 0 56028 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_609
timestamp 1
transform 1 0 57132 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_615
timestamp 1
transform 1 0 57684 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_617
timestamp 1636968456
transform 1 0 57868 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_629
timestamp 1636968456
transform 1 0 58972 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_641
timestamp 1636968456
transform 1 0 60076 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_653
timestamp 1636968456
transform 1 0 61180 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_665
timestamp 1
transform 1 0 62284 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_671
timestamp 1
transform 1 0 62836 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_673
timestamp 1636968456
transform 1 0 63020 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_685
timestamp 1636968456
transform 1 0 64124 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_697
timestamp 1636968456
transform 1 0 65228 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_709
timestamp 1636968456
transform 1 0 66332 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_721
timestamp 1
transform 1 0 67436 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_727
timestamp 1
transform 1 0 67988 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_729
timestamp 1636968456
transform 1 0 68172 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_741
timestamp 1636968456
transform 1 0 69276 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_753
timestamp 1636968456
transform 1 0 70380 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_765
timestamp 1636968456
transform 1 0 71484 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_777
timestamp 1
transform 1 0 72588 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_783
timestamp 1
transform 1 0 73140 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_785
timestamp 1636968456
transform 1 0 73324 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_797
timestamp 1636968456
transform 1 0 74428 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_809
timestamp 1636968456
transform 1 0 75532 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_821
timestamp 1636968456
transform 1 0 76636 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_833
timestamp 1
transform 1 0 77740 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_839
timestamp 1
transform 1 0 78292 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_841
timestamp 1636968456
transform 1 0 78476 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_853
timestamp 1636968456
transform 1 0 79580 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_865
timestamp 1636968456
transform 1 0 80684 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_877
timestamp 1636968456
transform 1 0 81788 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_889
timestamp 1
transform 1 0 82892 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_895
timestamp 1
transform 1 0 83444 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_897
timestamp 1636968456
transform 1 0 83628 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_909
timestamp 1636968456
transform 1 0 84732 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_921
timestamp 1636968456
transform 1 0 85836 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_933
timestamp 1636968456
transform 1 0 86940 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_945
timestamp 1
transform 1 0 88044 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_951
timestamp 1
transform 1 0 88596 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_953
timestamp 1636968456
transform 1 0 88780 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_965
timestamp 1636968456
transform 1 0 89884 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_977
timestamp 1636968456
transform 1 0 90988 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_989
timestamp 1636968456
transform 1 0 92092 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_1001
timestamp 1
transform 1 0 93196 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_1007
timestamp 1
transform 1 0 93748 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_1009
timestamp 1636968456
transform 1 0 93932 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_1021
timestamp 1636968456
transform 1 0 95036 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_1033
timestamp 1636968456
transform 1 0 96140 0 -1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_1045
timestamp 1636968456
transform 1 0 97244 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_121_1057
timestamp 1
transform 1 0 98348 0 -1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_121_1063
timestamp 1
transform 1 0 98900 0 -1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_1065
timestamp 1636968456
transform 1 0 99084 0 -1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_121_1077
timestamp 1
transform 1 0 100188 0 -1 68544
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_122_3
timestamp 1636968456
transform 1 0 1380 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_15
timestamp 1636968456
transform 1 0 2484 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_122_27
timestamp 1
transform 1 0 3588 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_29
timestamp 1636968456
transform 1 0 3772 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_41
timestamp 1636968456
transform 1 0 4876 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_53
timestamp 1636968456
transform 1 0 5980 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_65
timestamp 1636968456
transform 1 0 7084 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_77
timestamp 1
transform 1 0 8188 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_83
timestamp 1
transform 1 0 8740 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_85
timestamp 1636968456
transform 1 0 8924 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_97
timestamp 1636968456
transform 1 0 10028 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_109
timestamp 1636968456
transform 1 0 11132 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_121
timestamp 1636968456
transform 1 0 12236 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_133
timestamp 1
transform 1 0 13340 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_139
timestamp 1
transform 1 0 13892 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_141
timestamp 1636968456
transform 1 0 14076 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_153
timestamp 1636968456
transform 1 0 15180 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_165
timestamp 1636968456
transform 1 0 16284 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_177
timestamp 1636968456
transform 1 0 17388 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_189
timestamp 1
transform 1 0 18492 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_195
timestamp 1
transform 1 0 19044 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_197
timestamp 1636968456
transform 1 0 19228 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_209
timestamp 1636968456
transform 1 0 20332 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_221
timestamp 1636968456
transform 1 0 21436 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_233
timestamp 1636968456
transform 1 0 22540 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_245
timestamp 1
transform 1 0 23644 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_251
timestamp 1
transform 1 0 24196 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_253
timestamp 1636968456
transform 1 0 24380 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_265
timestamp 1636968456
transform 1 0 25484 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_277
timestamp 1636968456
transform 1 0 26588 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_289
timestamp 1636968456
transform 1 0 27692 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_301
timestamp 1
transform 1 0 28796 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_307
timestamp 1
transform 1 0 29348 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_309
timestamp 1636968456
transform 1 0 29532 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_321
timestamp 1636968456
transform 1 0 30636 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_333
timestamp 1636968456
transform 1 0 31740 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_345
timestamp 1636968456
transform 1 0 32844 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_357
timestamp 1
transform 1 0 33948 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_363
timestamp 1
transform 1 0 34500 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_365
timestamp 1636968456
transform 1 0 34684 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_377
timestamp 1636968456
transform 1 0 35788 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_389
timestamp 1636968456
transform 1 0 36892 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_401
timestamp 1636968456
transform 1 0 37996 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_413
timestamp 1
transform 1 0 39100 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_419
timestamp 1
transform 1 0 39652 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_421
timestamp 1636968456
transform 1 0 39836 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_433
timestamp 1636968456
transform 1 0 40940 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_445
timestamp 1636968456
transform 1 0 42044 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_457
timestamp 1636968456
transform 1 0 43148 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_469
timestamp 1
transform 1 0 44252 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_475
timestamp 1
transform 1 0 44804 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_477
timestamp 1636968456
transform 1 0 44988 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_489
timestamp 1636968456
transform 1 0 46092 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_501
timestamp 1636968456
transform 1 0 47196 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_513
timestamp 1636968456
transform 1 0 48300 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_525
timestamp 1
transform 1 0 49404 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_531
timestamp 1
transform 1 0 49956 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_533
timestamp 1636968456
transform 1 0 50140 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_545
timestamp 1636968456
transform 1 0 51244 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_557
timestamp 1636968456
transform 1 0 52348 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_569
timestamp 1636968456
transform 1 0 53452 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_581
timestamp 1
transform 1 0 54556 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_587
timestamp 1
transform 1 0 55108 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_589
timestamp 1636968456
transform 1 0 55292 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_601
timestamp 1636968456
transform 1 0 56396 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_613
timestamp 1636968456
transform 1 0 57500 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_625
timestamp 1636968456
transform 1 0 58604 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_637
timestamp 1
transform 1 0 59708 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_643
timestamp 1
transform 1 0 60260 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_645
timestamp 1636968456
transform 1 0 60444 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_657
timestamp 1636968456
transform 1 0 61548 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_669
timestamp 1636968456
transform 1 0 62652 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_681
timestamp 1636968456
transform 1 0 63756 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_693
timestamp 1
transform 1 0 64860 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_699
timestamp 1
transform 1 0 65412 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_701
timestamp 1636968456
transform 1 0 65596 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_713
timestamp 1636968456
transform 1 0 66700 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_725
timestamp 1636968456
transform 1 0 67804 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_737
timestamp 1636968456
transform 1 0 68908 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_749
timestamp 1
transform 1 0 70012 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_755
timestamp 1
transform 1 0 70564 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_757
timestamp 1636968456
transform 1 0 70748 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_769
timestamp 1636968456
transform 1 0 71852 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_781
timestamp 1636968456
transform 1 0 72956 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_793
timestamp 1636968456
transform 1 0 74060 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_805
timestamp 1
transform 1 0 75164 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_811
timestamp 1
transform 1 0 75716 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_813
timestamp 1636968456
transform 1 0 75900 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_825
timestamp 1636968456
transform 1 0 77004 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_837
timestamp 1636968456
transform 1 0 78108 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_849
timestamp 1636968456
transform 1 0 79212 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_861
timestamp 1
transform 1 0 80316 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_867
timestamp 1
transform 1 0 80868 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_869
timestamp 1636968456
transform 1 0 81052 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_881
timestamp 1636968456
transform 1 0 82156 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_893
timestamp 1636968456
transform 1 0 83260 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_905
timestamp 1636968456
transform 1 0 84364 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_917
timestamp 1
transform 1 0 85468 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_923
timestamp 1
transform 1 0 86020 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_925
timestamp 1636968456
transform 1 0 86204 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_937
timestamp 1636968456
transform 1 0 87308 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_949
timestamp 1636968456
transform 1 0 88412 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_961
timestamp 1636968456
transform 1 0 89516 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_973
timestamp 1
transform 1 0 90620 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_979
timestamp 1
transform 1 0 91172 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_981
timestamp 1636968456
transform 1 0 91356 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_993
timestamp 1636968456
transform 1 0 92460 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_1005
timestamp 1636968456
transform 1 0 93564 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_1017
timestamp 1636968456
transform 1 0 94668 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_1029
timestamp 1
transform 1 0 95772 0 1 68544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_122_1035
timestamp 1
transform 1 0 96324 0 1 68544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_1037
timestamp 1636968456
transform 1 0 96508 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_1049
timestamp 1636968456
transform 1 0 97612 0 1 68544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_1061
timestamp 1636968456
transform 1 0 98716 0 1 68544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_122_1073
timestamp 1
transform 1 0 99820 0 1 68544
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_123_3
timestamp 1636968456
transform 1 0 1380 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_15
timestamp 1636968456
transform 1 0 2484 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_27
timestamp 1636968456
transform 1 0 3588 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_39
timestamp 1636968456
transform 1 0 4692 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_123_51
timestamp 1
transform 1 0 5796 0 -1 69632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_123_55
timestamp 1
transform 1 0 6164 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_57
timestamp 1636968456
transform 1 0 6348 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_69
timestamp 1636968456
transform 1 0 7452 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_81
timestamp 1636968456
transform 1 0 8556 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_93
timestamp 1636968456
transform 1 0 9660 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_105
timestamp 1
transform 1 0 10764 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_111
timestamp 1
transform 1 0 11316 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_113
timestamp 1636968456
transform 1 0 11500 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_125
timestamp 1636968456
transform 1 0 12604 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_137
timestamp 1636968456
transform 1 0 13708 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_149
timestamp 1636968456
transform 1 0 14812 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_161
timestamp 1
transform 1 0 15916 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_167
timestamp 1
transform 1 0 16468 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_169
timestamp 1636968456
transform 1 0 16652 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_181
timestamp 1636968456
transform 1 0 17756 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_193
timestamp 1636968456
transform 1 0 18860 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_205
timestamp 1636968456
transform 1 0 19964 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_217
timestamp 1
transform 1 0 21068 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_223
timestamp 1
transform 1 0 21620 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_225
timestamp 1636968456
transform 1 0 21804 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_237
timestamp 1636968456
transform 1 0 22908 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_249
timestamp 1636968456
transform 1 0 24012 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_261
timestamp 1636968456
transform 1 0 25116 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_273
timestamp 1
transform 1 0 26220 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_279
timestamp 1
transform 1 0 26772 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_281
timestamp 1636968456
transform 1 0 26956 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_293
timestamp 1636968456
transform 1 0 28060 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_305
timestamp 1636968456
transform 1 0 29164 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_317
timestamp 1636968456
transform 1 0 30268 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_329
timestamp 1
transform 1 0 31372 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_335
timestamp 1
transform 1 0 31924 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_337
timestamp 1636968456
transform 1 0 32108 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_349
timestamp 1636968456
transform 1 0 33212 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_361
timestamp 1636968456
transform 1 0 34316 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_373
timestamp 1636968456
transform 1 0 35420 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_385
timestamp 1
transform 1 0 36524 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_391
timestamp 1
transform 1 0 37076 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_393
timestamp 1636968456
transform 1 0 37260 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_405
timestamp 1636968456
transform 1 0 38364 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_417
timestamp 1636968456
transform 1 0 39468 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_429
timestamp 1636968456
transform 1 0 40572 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_441
timestamp 1
transform 1 0 41676 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_447
timestamp 1
transform 1 0 42228 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_449
timestamp 1636968456
transform 1 0 42412 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_461
timestamp 1636968456
transform 1 0 43516 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_473
timestamp 1636968456
transform 1 0 44620 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_485
timestamp 1636968456
transform 1 0 45724 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_497
timestamp 1
transform 1 0 46828 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_503
timestamp 1
transform 1 0 47380 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_505
timestamp 1636968456
transform 1 0 47564 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_517
timestamp 1636968456
transform 1 0 48668 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_529
timestamp 1636968456
transform 1 0 49772 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_541
timestamp 1636968456
transform 1 0 50876 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_553
timestamp 1
transform 1 0 51980 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_559
timestamp 1
transform 1 0 52532 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_561
timestamp 1636968456
transform 1 0 52716 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_573
timestamp 1636968456
transform 1 0 53820 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_585
timestamp 1636968456
transform 1 0 54924 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_597
timestamp 1636968456
transform 1 0 56028 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_609
timestamp 1
transform 1 0 57132 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_615
timestamp 1
transform 1 0 57684 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_617
timestamp 1636968456
transform 1 0 57868 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_629
timestamp 1636968456
transform 1 0 58972 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_641
timestamp 1636968456
transform 1 0 60076 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_653
timestamp 1636968456
transform 1 0 61180 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_665
timestamp 1
transform 1 0 62284 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_671
timestamp 1
transform 1 0 62836 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_673
timestamp 1636968456
transform 1 0 63020 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_685
timestamp 1636968456
transform 1 0 64124 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_697
timestamp 1636968456
transform 1 0 65228 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_709
timestamp 1636968456
transform 1 0 66332 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_721
timestamp 1
transform 1 0 67436 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_727
timestamp 1
transform 1 0 67988 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_729
timestamp 1636968456
transform 1 0 68172 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_741
timestamp 1636968456
transform 1 0 69276 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_753
timestamp 1636968456
transform 1 0 70380 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_765
timestamp 1636968456
transform 1 0 71484 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_777
timestamp 1
transform 1 0 72588 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_783
timestamp 1
transform 1 0 73140 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_785
timestamp 1636968456
transform 1 0 73324 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_797
timestamp 1636968456
transform 1 0 74428 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_809
timestamp 1636968456
transform 1 0 75532 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_821
timestamp 1636968456
transform 1 0 76636 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_833
timestamp 1
transform 1 0 77740 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_839
timestamp 1
transform 1 0 78292 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_841
timestamp 1636968456
transform 1 0 78476 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_853
timestamp 1636968456
transform 1 0 79580 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_865
timestamp 1636968456
transform 1 0 80684 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_877
timestamp 1636968456
transform 1 0 81788 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_889
timestamp 1
transform 1 0 82892 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_895
timestamp 1
transform 1 0 83444 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_897
timestamp 1636968456
transform 1 0 83628 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_909
timestamp 1636968456
transform 1 0 84732 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_921
timestamp 1636968456
transform 1 0 85836 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_933
timestamp 1636968456
transform 1 0 86940 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_945
timestamp 1
transform 1 0 88044 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_951
timestamp 1
transform 1 0 88596 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_953
timestamp 1636968456
transform 1 0 88780 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_965
timestamp 1636968456
transform 1 0 89884 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_977
timestamp 1636968456
transform 1 0 90988 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_989
timestamp 1636968456
transform 1 0 92092 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_1001
timestamp 1
transform 1 0 93196 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_1007
timestamp 1
transform 1 0 93748 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_1009
timestamp 1636968456
transform 1 0 93932 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_1021
timestamp 1636968456
transform 1 0 95036 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_1033
timestamp 1636968456
transform 1 0 96140 0 -1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_123_1045
timestamp 1636968456
transform 1 0 97244 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_123_1057
timestamp 1
transform 1 0 98348 0 -1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_123_1063
timestamp 1
transform 1 0 98900 0 -1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_1065
timestamp 1636968456
transform 1 0 99084 0 -1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_123_1077
timestamp 1
transform 1 0 100188 0 -1 69632
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_124_3
timestamp 1636968456
transform 1 0 1380 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_15
timestamp 1636968456
transform 1 0 2484 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_124_27
timestamp 1
transform 1 0 3588 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_29
timestamp 1636968456
transform 1 0 3772 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_41
timestamp 1636968456
transform 1 0 4876 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_53
timestamp 1636968456
transform 1 0 5980 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_65
timestamp 1636968456
transform 1 0 7084 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_77
timestamp 1
transform 1 0 8188 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_83
timestamp 1
transform 1 0 8740 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_85
timestamp 1636968456
transform 1 0 8924 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_97
timestamp 1636968456
transform 1 0 10028 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_109
timestamp 1636968456
transform 1 0 11132 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_121
timestamp 1636968456
transform 1 0 12236 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_133
timestamp 1
transform 1 0 13340 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_139
timestamp 1
transform 1 0 13892 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_141
timestamp 1636968456
transform 1 0 14076 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_153
timestamp 1636968456
transform 1 0 15180 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_165
timestamp 1636968456
transform 1 0 16284 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_177
timestamp 1636968456
transform 1 0 17388 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_189
timestamp 1
transform 1 0 18492 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_195
timestamp 1
transform 1 0 19044 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_197
timestamp 1636968456
transform 1 0 19228 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_209
timestamp 1636968456
transform 1 0 20332 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_221
timestamp 1636968456
transform 1 0 21436 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_233
timestamp 1636968456
transform 1 0 22540 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_245
timestamp 1
transform 1 0 23644 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_251
timestamp 1
transform 1 0 24196 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_253
timestamp 1636968456
transform 1 0 24380 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_265
timestamp 1636968456
transform 1 0 25484 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_277
timestamp 1636968456
transform 1 0 26588 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_289
timestamp 1636968456
transform 1 0 27692 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_301
timestamp 1
transform 1 0 28796 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_307
timestamp 1
transform 1 0 29348 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_309
timestamp 1636968456
transform 1 0 29532 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_321
timestamp 1636968456
transform 1 0 30636 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_333
timestamp 1636968456
transform 1 0 31740 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_345
timestamp 1636968456
transform 1 0 32844 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_357
timestamp 1
transform 1 0 33948 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_363
timestamp 1
transform 1 0 34500 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_365
timestamp 1636968456
transform 1 0 34684 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_377
timestamp 1636968456
transform 1 0 35788 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_389
timestamp 1636968456
transform 1 0 36892 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_401
timestamp 1636968456
transform 1 0 37996 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_413
timestamp 1
transform 1 0 39100 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_419
timestamp 1
transform 1 0 39652 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_421
timestamp 1636968456
transform 1 0 39836 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_433
timestamp 1636968456
transform 1 0 40940 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_445
timestamp 1636968456
transform 1 0 42044 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_457
timestamp 1636968456
transform 1 0 43148 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_469
timestamp 1
transform 1 0 44252 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_475
timestamp 1
transform 1 0 44804 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_477
timestamp 1636968456
transform 1 0 44988 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_489
timestamp 1636968456
transform 1 0 46092 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_501
timestamp 1636968456
transform 1 0 47196 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_513
timestamp 1636968456
transform 1 0 48300 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_525
timestamp 1
transform 1 0 49404 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_531
timestamp 1
transform 1 0 49956 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_533
timestamp 1636968456
transform 1 0 50140 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_545
timestamp 1636968456
transform 1 0 51244 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_557
timestamp 1636968456
transform 1 0 52348 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_569
timestamp 1636968456
transform 1 0 53452 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_581
timestamp 1
transform 1 0 54556 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_587
timestamp 1
transform 1 0 55108 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_589
timestamp 1636968456
transform 1 0 55292 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_601
timestamp 1636968456
transform 1 0 56396 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_613
timestamp 1636968456
transform 1 0 57500 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_625
timestamp 1636968456
transform 1 0 58604 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_637
timestamp 1
transform 1 0 59708 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_643
timestamp 1
transform 1 0 60260 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_645
timestamp 1636968456
transform 1 0 60444 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_657
timestamp 1636968456
transform 1 0 61548 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_669
timestamp 1636968456
transform 1 0 62652 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_681
timestamp 1636968456
transform 1 0 63756 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_693
timestamp 1
transform 1 0 64860 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_699
timestamp 1
transform 1 0 65412 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_701
timestamp 1636968456
transform 1 0 65596 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_713
timestamp 1636968456
transform 1 0 66700 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_725
timestamp 1636968456
transform 1 0 67804 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_737
timestamp 1636968456
transform 1 0 68908 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_749
timestamp 1
transform 1 0 70012 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_755
timestamp 1
transform 1 0 70564 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_757
timestamp 1636968456
transform 1 0 70748 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_769
timestamp 1636968456
transform 1 0 71852 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_781
timestamp 1636968456
transform 1 0 72956 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_793
timestamp 1636968456
transform 1 0 74060 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_805
timestamp 1
transform 1 0 75164 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_811
timestamp 1
transform 1 0 75716 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_813
timestamp 1636968456
transform 1 0 75900 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_825
timestamp 1636968456
transform 1 0 77004 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_837
timestamp 1636968456
transform 1 0 78108 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_849
timestamp 1636968456
transform 1 0 79212 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_861
timestamp 1
transform 1 0 80316 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_867
timestamp 1
transform 1 0 80868 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_869
timestamp 1636968456
transform 1 0 81052 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_881
timestamp 1636968456
transform 1 0 82156 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_893
timestamp 1636968456
transform 1 0 83260 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_905
timestamp 1636968456
transform 1 0 84364 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_917
timestamp 1
transform 1 0 85468 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_923
timestamp 1
transform 1 0 86020 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_925
timestamp 1636968456
transform 1 0 86204 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_937
timestamp 1636968456
transform 1 0 87308 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_949
timestamp 1636968456
transform 1 0 88412 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_961
timestamp 1636968456
transform 1 0 89516 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_973
timestamp 1
transform 1 0 90620 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_979
timestamp 1
transform 1 0 91172 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_981
timestamp 1636968456
transform 1 0 91356 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_993
timestamp 1636968456
transform 1 0 92460 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_1005
timestamp 1636968456
transform 1 0 93564 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_1017
timestamp 1636968456
transform 1 0 94668 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_124_1029
timestamp 1
transform 1 0 95772 0 1 69632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_124_1035
timestamp 1
transform 1 0 96324 0 1 69632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_1037
timestamp 1636968456
transform 1 0 96508 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_1049
timestamp 1636968456
transform 1 0 97612 0 1 69632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_1061
timestamp 1636968456
transform 1 0 98716 0 1 69632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_124_1073
timestamp 1
transform 1 0 99820 0 1 69632
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_125_3
timestamp 1636968456
transform 1 0 1380 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_15
timestamp 1636968456
transform 1 0 2484 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_27
timestamp 1636968456
transform 1 0 3588 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_39
timestamp 1636968456
transform 1 0 4692 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_125_51
timestamp 1
transform 1 0 5796 0 -1 70720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_125_55
timestamp 1
transform 1 0 6164 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_57
timestamp 1636968456
transform 1 0 6348 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_69
timestamp 1636968456
transform 1 0 7452 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_81
timestamp 1636968456
transform 1 0 8556 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_93
timestamp 1636968456
transform 1 0 9660 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_105
timestamp 1
transform 1 0 10764 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_111
timestamp 1
transform 1 0 11316 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_113
timestamp 1636968456
transform 1 0 11500 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_125
timestamp 1636968456
transform 1 0 12604 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_137
timestamp 1636968456
transform 1 0 13708 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_149
timestamp 1636968456
transform 1 0 14812 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_161
timestamp 1
transform 1 0 15916 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_167
timestamp 1
transform 1 0 16468 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_169
timestamp 1636968456
transform 1 0 16652 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_181
timestamp 1636968456
transform 1 0 17756 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_193
timestamp 1636968456
transform 1 0 18860 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_205
timestamp 1636968456
transform 1 0 19964 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_217
timestamp 1
transform 1 0 21068 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_223
timestamp 1
transform 1 0 21620 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_225
timestamp 1636968456
transform 1 0 21804 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_237
timestamp 1636968456
transform 1 0 22908 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_249
timestamp 1636968456
transform 1 0 24012 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_261
timestamp 1636968456
transform 1 0 25116 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_273
timestamp 1
transform 1 0 26220 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_279
timestamp 1
transform 1 0 26772 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_281
timestamp 1636968456
transform 1 0 26956 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_293
timestamp 1636968456
transform 1 0 28060 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_305
timestamp 1636968456
transform 1 0 29164 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_317
timestamp 1636968456
transform 1 0 30268 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_329
timestamp 1
transform 1 0 31372 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_335
timestamp 1
transform 1 0 31924 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_337
timestamp 1636968456
transform 1 0 32108 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_349
timestamp 1636968456
transform 1 0 33212 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_361
timestamp 1636968456
transform 1 0 34316 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_373
timestamp 1636968456
transform 1 0 35420 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_385
timestamp 1
transform 1 0 36524 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_391
timestamp 1
transform 1 0 37076 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_393
timestamp 1636968456
transform 1 0 37260 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_405
timestamp 1636968456
transform 1 0 38364 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_417
timestamp 1636968456
transform 1 0 39468 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_429
timestamp 1636968456
transform 1 0 40572 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_441
timestamp 1
transform 1 0 41676 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_447
timestamp 1
transform 1 0 42228 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_449
timestamp 1636968456
transform 1 0 42412 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_461
timestamp 1636968456
transform 1 0 43516 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_473
timestamp 1636968456
transform 1 0 44620 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_485
timestamp 1636968456
transform 1 0 45724 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_497
timestamp 1
transform 1 0 46828 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_503
timestamp 1
transform 1 0 47380 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_505
timestamp 1636968456
transform 1 0 47564 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_517
timestamp 1636968456
transform 1 0 48668 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_529
timestamp 1636968456
transform 1 0 49772 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_541
timestamp 1636968456
transform 1 0 50876 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_553
timestamp 1
transform 1 0 51980 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_559
timestamp 1
transform 1 0 52532 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_561
timestamp 1636968456
transform 1 0 52716 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_573
timestamp 1636968456
transform 1 0 53820 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_585
timestamp 1636968456
transform 1 0 54924 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_597
timestamp 1636968456
transform 1 0 56028 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_609
timestamp 1
transform 1 0 57132 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_615
timestamp 1
transform 1 0 57684 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_617
timestamp 1636968456
transform 1 0 57868 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_629
timestamp 1636968456
transform 1 0 58972 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_641
timestamp 1636968456
transform 1 0 60076 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_653
timestamp 1636968456
transform 1 0 61180 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_665
timestamp 1
transform 1 0 62284 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_671
timestamp 1
transform 1 0 62836 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_673
timestamp 1636968456
transform 1 0 63020 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_685
timestamp 1636968456
transform 1 0 64124 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_697
timestamp 1636968456
transform 1 0 65228 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_709
timestamp 1636968456
transform 1 0 66332 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_721
timestamp 1
transform 1 0 67436 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_727
timestamp 1
transform 1 0 67988 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_729
timestamp 1636968456
transform 1 0 68172 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_741
timestamp 1636968456
transform 1 0 69276 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_753
timestamp 1636968456
transform 1 0 70380 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_765
timestamp 1636968456
transform 1 0 71484 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_777
timestamp 1
transform 1 0 72588 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_783
timestamp 1
transform 1 0 73140 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_785
timestamp 1636968456
transform 1 0 73324 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_797
timestamp 1636968456
transform 1 0 74428 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_809
timestamp 1636968456
transform 1 0 75532 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_821
timestamp 1636968456
transform 1 0 76636 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_833
timestamp 1
transform 1 0 77740 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_839
timestamp 1
transform 1 0 78292 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_841
timestamp 1636968456
transform 1 0 78476 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_853
timestamp 1636968456
transform 1 0 79580 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_865
timestamp 1636968456
transform 1 0 80684 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_877
timestamp 1636968456
transform 1 0 81788 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_889
timestamp 1
transform 1 0 82892 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_895
timestamp 1
transform 1 0 83444 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_897
timestamp 1636968456
transform 1 0 83628 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_909
timestamp 1636968456
transform 1 0 84732 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_921
timestamp 1636968456
transform 1 0 85836 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_933
timestamp 1636968456
transform 1 0 86940 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_945
timestamp 1
transform 1 0 88044 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_951
timestamp 1
transform 1 0 88596 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_953
timestamp 1636968456
transform 1 0 88780 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_965
timestamp 1636968456
transform 1 0 89884 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_977
timestamp 1636968456
transform 1 0 90988 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_989
timestamp 1636968456
transform 1 0 92092 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_1001
timestamp 1
transform 1 0 93196 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_1007
timestamp 1
transform 1 0 93748 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_1009
timestamp 1636968456
transform 1 0 93932 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_1021
timestamp 1636968456
transform 1 0 95036 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_1033
timestamp 1636968456
transform 1 0 96140 0 -1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_125_1045
timestamp 1636968456
transform 1 0 97244 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_125_1057
timestamp 1
transform 1 0 98348 0 -1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_125_1063
timestamp 1
transform 1 0 98900 0 -1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_1065
timestamp 1636968456
transform 1 0 99084 0 -1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_125_1077
timestamp 1
transform 1 0 100188 0 -1 70720
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_126_3
timestamp 1636968456
transform 1 0 1380 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_15
timestamp 1636968456
transform 1 0 2484 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_126_27
timestamp 1
transform 1 0 3588 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_29
timestamp 1636968456
transform 1 0 3772 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_41
timestamp 1636968456
transform 1 0 4876 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_53
timestamp 1636968456
transform 1 0 5980 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_65
timestamp 1636968456
transform 1 0 7084 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_77
timestamp 1
transform 1 0 8188 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_83
timestamp 1
transform 1 0 8740 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_85
timestamp 1636968456
transform 1 0 8924 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_97
timestamp 1636968456
transform 1 0 10028 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_109
timestamp 1636968456
transform 1 0 11132 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_121
timestamp 1636968456
transform 1 0 12236 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_133
timestamp 1
transform 1 0 13340 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_139
timestamp 1
transform 1 0 13892 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_141
timestamp 1636968456
transform 1 0 14076 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_153
timestamp 1636968456
transform 1 0 15180 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_165
timestamp 1636968456
transform 1 0 16284 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_177
timestamp 1636968456
transform 1 0 17388 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_189
timestamp 1
transform 1 0 18492 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_195
timestamp 1
transform 1 0 19044 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_197
timestamp 1636968456
transform 1 0 19228 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_209
timestamp 1636968456
transform 1 0 20332 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_221
timestamp 1636968456
transform 1 0 21436 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_233
timestamp 1636968456
transform 1 0 22540 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_245
timestamp 1
transform 1 0 23644 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_251
timestamp 1
transform 1 0 24196 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_253
timestamp 1636968456
transform 1 0 24380 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_265
timestamp 1636968456
transform 1 0 25484 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_277
timestamp 1636968456
transform 1 0 26588 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_289
timestamp 1636968456
transform 1 0 27692 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_301
timestamp 1
transform 1 0 28796 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_307
timestamp 1
transform 1 0 29348 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_309
timestamp 1636968456
transform 1 0 29532 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_321
timestamp 1636968456
transform 1 0 30636 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_333
timestamp 1636968456
transform 1 0 31740 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_345
timestamp 1636968456
transform 1 0 32844 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_357
timestamp 1
transform 1 0 33948 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_363
timestamp 1
transform 1 0 34500 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_365
timestamp 1636968456
transform 1 0 34684 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_377
timestamp 1636968456
transform 1 0 35788 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_389
timestamp 1636968456
transform 1 0 36892 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_401
timestamp 1636968456
transform 1 0 37996 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_413
timestamp 1
transform 1 0 39100 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_419
timestamp 1
transform 1 0 39652 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_421
timestamp 1636968456
transform 1 0 39836 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_433
timestamp 1636968456
transform 1 0 40940 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_445
timestamp 1636968456
transform 1 0 42044 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_457
timestamp 1636968456
transform 1 0 43148 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_469
timestamp 1
transform 1 0 44252 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_475
timestamp 1
transform 1 0 44804 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_477
timestamp 1636968456
transform 1 0 44988 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_489
timestamp 1636968456
transform 1 0 46092 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_501
timestamp 1636968456
transform 1 0 47196 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_513
timestamp 1636968456
transform 1 0 48300 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_525
timestamp 1
transform 1 0 49404 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_531
timestamp 1
transform 1 0 49956 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_533
timestamp 1636968456
transform 1 0 50140 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_545
timestamp 1636968456
transform 1 0 51244 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_557
timestamp 1636968456
transform 1 0 52348 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_569
timestamp 1636968456
transform 1 0 53452 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_581
timestamp 1
transform 1 0 54556 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_587
timestamp 1
transform 1 0 55108 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_589
timestamp 1636968456
transform 1 0 55292 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_601
timestamp 1636968456
transform 1 0 56396 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_613
timestamp 1636968456
transform 1 0 57500 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_625
timestamp 1636968456
transform 1 0 58604 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_637
timestamp 1
transform 1 0 59708 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_643
timestamp 1
transform 1 0 60260 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_645
timestamp 1636968456
transform 1 0 60444 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_657
timestamp 1636968456
transform 1 0 61548 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_669
timestamp 1636968456
transform 1 0 62652 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_681
timestamp 1636968456
transform 1 0 63756 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_693
timestamp 1
transform 1 0 64860 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_699
timestamp 1
transform 1 0 65412 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_701
timestamp 1636968456
transform 1 0 65596 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_713
timestamp 1636968456
transform 1 0 66700 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_725
timestamp 1636968456
transform 1 0 67804 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_737
timestamp 1636968456
transform 1 0 68908 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_749
timestamp 1
transform 1 0 70012 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_755
timestamp 1
transform 1 0 70564 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_757
timestamp 1636968456
transform 1 0 70748 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_769
timestamp 1636968456
transform 1 0 71852 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_781
timestamp 1636968456
transform 1 0 72956 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_793
timestamp 1636968456
transform 1 0 74060 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_805
timestamp 1
transform 1 0 75164 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_811
timestamp 1
transform 1 0 75716 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_813
timestamp 1636968456
transform 1 0 75900 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_825
timestamp 1636968456
transform 1 0 77004 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_837
timestamp 1636968456
transform 1 0 78108 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_849
timestamp 1636968456
transform 1 0 79212 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_861
timestamp 1
transform 1 0 80316 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_867
timestamp 1
transform 1 0 80868 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_869
timestamp 1636968456
transform 1 0 81052 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_881
timestamp 1636968456
transform 1 0 82156 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_893
timestamp 1636968456
transform 1 0 83260 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_905
timestamp 1636968456
transform 1 0 84364 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_917
timestamp 1
transform 1 0 85468 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_923
timestamp 1
transform 1 0 86020 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_925
timestamp 1636968456
transform 1 0 86204 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_937
timestamp 1636968456
transform 1 0 87308 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_949
timestamp 1636968456
transform 1 0 88412 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_961
timestamp 1636968456
transform 1 0 89516 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_973
timestamp 1
transform 1 0 90620 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_979
timestamp 1
transform 1 0 91172 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_981
timestamp 1636968456
transform 1 0 91356 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_993
timestamp 1636968456
transform 1 0 92460 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_1005
timestamp 1636968456
transform 1 0 93564 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_1017
timestamp 1636968456
transform 1 0 94668 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_1029
timestamp 1
transform 1 0 95772 0 1 70720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_126_1035
timestamp 1
transform 1 0 96324 0 1 70720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_1037
timestamp 1636968456
transform 1 0 96508 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_1049
timestamp 1636968456
transform 1 0 97612 0 1 70720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_1061
timestamp 1636968456
transform 1 0 98716 0 1 70720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_126_1073
timestamp 1
transform 1 0 99820 0 1 70720
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_127_3
timestamp 1636968456
transform 1 0 1380 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_15
timestamp 1636968456
transform 1 0 2484 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_27
timestamp 1636968456
transform 1 0 3588 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_39
timestamp 1636968456
transform 1 0 4692 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_127_51
timestamp 1
transform 1 0 5796 0 -1 71808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_127_55
timestamp 1
transform 1 0 6164 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_57
timestamp 1636968456
transform 1 0 6348 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_69
timestamp 1636968456
transform 1 0 7452 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_81
timestamp 1636968456
transform 1 0 8556 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_93
timestamp 1636968456
transform 1 0 9660 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_105
timestamp 1
transform 1 0 10764 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_111
timestamp 1
transform 1 0 11316 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_113
timestamp 1636968456
transform 1 0 11500 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_125
timestamp 1636968456
transform 1 0 12604 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_137
timestamp 1636968456
transform 1 0 13708 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_149
timestamp 1636968456
transform 1 0 14812 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_161
timestamp 1
transform 1 0 15916 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_167
timestamp 1
transform 1 0 16468 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_169
timestamp 1636968456
transform 1 0 16652 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_181
timestamp 1636968456
transform 1 0 17756 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_193
timestamp 1636968456
transform 1 0 18860 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_205
timestamp 1636968456
transform 1 0 19964 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_217
timestamp 1
transform 1 0 21068 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_223
timestamp 1
transform 1 0 21620 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_225
timestamp 1636968456
transform 1 0 21804 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_237
timestamp 1636968456
transform 1 0 22908 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_249
timestamp 1636968456
transform 1 0 24012 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_261
timestamp 1636968456
transform 1 0 25116 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_273
timestamp 1
transform 1 0 26220 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_279
timestamp 1
transform 1 0 26772 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_281
timestamp 1636968456
transform 1 0 26956 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_293
timestamp 1636968456
transform 1 0 28060 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_305
timestamp 1636968456
transform 1 0 29164 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_317
timestamp 1636968456
transform 1 0 30268 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_329
timestamp 1
transform 1 0 31372 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_335
timestamp 1
transform 1 0 31924 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_337
timestamp 1636968456
transform 1 0 32108 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_349
timestamp 1636968456
transform 1 0 33212 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_361
timestamp 1636968456
transform 1 0 34316 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_373
timestamp 1636968456
transform 1 0 35420 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_385
timestamp 1
transform 1 0 36524 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_391
timestamp 1
transform 1 0 37076 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_393
timestamp 1636968456
transform 1 0 37260 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_405
timestamp 1636968456
transform 1 0 38364 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_417
timestamp 1636968456
transform 1 0 39468 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_429
timestamp 1636968456
transform 1 0 40572 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_441
timestamp 1
transform 1 0 41676 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_447
timestamp 1
transform 1 0 42228 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_449
timestamp 1636968456
transform 1 0 42412 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_461
timestamp 1636968456
transform 1 0 43516 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_473
timestamp 1636968456
transform 1 0 44620 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_485
timestamp 1636968456
transform 1 0 45724 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_497
timestamp 1
transform 1 0 46828 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_503
timestamp 1
transform 1 0 47380 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_505
timestamp 1636968456
transform 1 0 47564 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_517
timestamp 1636968456
transform 1 0 48668 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_529
timestamp 1636968456
transform 1 0 49772 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_541
timestamp 1636968456
transform 1 0 50876 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_553
timestamp 1
transform 1 0 51980 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_559
timestamp 1
transform 1 0 52532 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_561
timestamp 1636968456
transform 1 0 52716 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_573
timestamp 1636968456
transform 1 0 53820 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_585
timestamp 1636968456
transform 1 0 54924 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_597
timestamp 1636968456
transform 1 0 56028 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_609
timestamp 1
transform 1 0 57132 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_615
timestamp 1
transform 1 0 57684 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_617
timestamp 1636968456
transform 1 0 57868 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_629
timestamp 1636968456
transform 1 0 58972 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_641
timestamp 1636968456
transform 1 0 60076 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_653
timestamp 1636968456
transform 1 0 61180 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_665
timestamp 1
transform 1 0 62284 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_671
timestamp 1
transform 1 0 62836 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_673
timestamp 1636968456
transform 1 0 63020 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_685
timestamp 1636968456
transform 1 0 64124 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_697
timestamp 1636968456
transform 1 0 65228 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_709
timestamp 1636968456
transform 1 0 66332 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_721
timestamp 1
transform 1 0 67436 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_727
timestamp 1
transform 1 0 67988 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_729
timestamp 1636968456
transform 1 0 68172 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_741
timestamp 1636968456
transform 1 0 69276 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_753
timestamp 1636968456
transform 1 0 70380 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_765
timestamp 1636968456
transform 1 0 71484 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_777
timestamp 1
transform 1 0 72588 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_783
timestamp 1
transform 1 0 73140 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_785
timestamp 1636968456
transform 1 0 73324 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_797
timestamp 1636968456
transform 1 0 74428 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_809
timestamp 1636968456
transform 1 0 75532 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_821
timestamp 1636968456
transform 1 0 76636 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_833
timestamp 1
transform 1 0 77740 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_839
timestamp 1
transform 1 0 78292 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_841
timestamp 1636968456
transform 1 0 78476 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_853
timestamp 1636968456
transform 1 0 79580 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_865
timestamp 1636968456
transform 1 0 80684 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_877
timestamp 1636968456
transform 1 0 81788 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_889
timestamp 1
transform 1 0 82892 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_895
timestamp 1
transform 1 0 83444 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_897
timestamp 1636968456
transform 1 0 83628 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_909
timestamp 1636968456
transform 1 0 84732 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_921
timestamp 1636968456
transform 1 0 85836 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_933
timestamp 1636968456
transform 1 0 86940 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_945
timestamp 1
transform 1 0 88044 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_951
timestamp 1
transform 1 0 88596 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_953
timestamp 1636968456
transform 1 0 88780 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_965
timestamp 1636968456
transform 1 0 89884 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_977
timestamp 1636968456
transform 1 0 90988 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_989
timestamp 1636968456
transform 1 0 92092 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_1001
timestamp 1
transform 1 0 93196 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_1007
timestamp 1
transform 1 0 93748 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_1009
timestamp 1636968456
transform 1 0 93932 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_1021
timestamp 1636968456
transform 1 0 95036 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_1033
timestamp 1636968456
transform 1 0 96140 0 -1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_127_1045
timestamp 1636968456
transform 1 0 97244 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_127_1057
timestamp 1
transform 1 0 98348 0 -1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_127_1063
timestamp 1
transform 1 0 98900 0 -1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_1065
timestamp 1636968456
transform 1 0 99084 0 -1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_127_1077
timestamp 1
transform 1 0 100188 0 -1 71808
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_128_3
timestamp 1636968456
transform 1 0 1380 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_15
timestamp 1636968456
transform 1 0 2484 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_128_27
timestamp 1
transform 1 0 3588 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_29
timestamp 1636968456
transform 1 0 3772 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_41
timestamp 1636968456
transform 1 0 4876 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_53
timestamp 1636968456
transform 1 0 5980 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_65
timestamp 1636968456
transform 1 0 7084 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_77
timestamp 1
transform 1 0 8188 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_83
timestamp 1
transform 1 0 8740 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_85
timestamp 1636968456
transform 1 0 8924 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_97
timestamp 1636968456
transform 1 0 10028 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_109
timestamp 1636968456
transform 1 0 11132 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_121
timestamp 1636968456
transform 1 0 12236 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_133
timestamp 1
transform 1 0 13340 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_139
timestamp 1
transform 1 0 13892 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_141
timestamp 1636968456
transform 1 0 14076 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_153
timestamp 1636968456
transform 1 0 15180 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_165
timestamp 1636968456
transform 1 0 16284 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_177
timestamp 1636968456
transform 1 0 17388 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_189
timestamp 1
transform 1 0 18492 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_195
timestamp 1
transform 1 0 19044 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_197
timestamp 1636968456
transform 1 0 19228 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_209
timestamp 1636968456
transform 1 0 20332 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_221
timestamp 1636968456
transform 1 0 21436 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_233
timestamp 1636968456
transform 1 0 22540 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_245
timestamp 1
transform 1 0 23644 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_251
timestamp 1
transform 1 0 24196 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_253
timestamp 1636968456
transform 1 0 24380 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_265
timestamp 1636968456
transform 1 0 25484 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_277
timestamp 1636968456
transform 1 0 26588 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_289
timestamp 1636968456
transform 1 0 27692 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_301
timestamp 1
transform 1 0 28796 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_307
timestamp 1
transform 1 0 29348 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_309
timestamp 1636968456
transform 1 0 29532 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_321
timestamp 1636968456
transform 1 0 30636 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_333
timestamp 1636968456
transform 1 0 31740 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_345
timestamp 1636968456
transform 1 0 32844 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_357
timestamp 1
transform 1 0 33948 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_363
timestamp 1
transform 1 0 34500 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_365
timestamp 1636968456
transform 1 0 34684 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_377
timestamp 1636968456
transform 1 0 35788 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_389
timestamp 1636968456
transform 1 0 36892 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_401
timestamp 1636968456
transform 1 0 37996 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_413
timestamp 1
transform 1 0 39100 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_419
timestamp 1
transform 1 0 39652 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_421
timestamp 1636968456
transform 1 0 39836 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_433
timestamp 1636968456
transform 1 0 40940 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_445
timestamp 1636968456
transform 1 0 42044 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_457
timestamp 1636968456
transform 1 0 43148 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_469
timestamp 1
transform 1 0 44252 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_475
timestamp 1
transform 1 0 44804 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_477
timestamp 1636968456
transform 1 0 44988 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_489
timestamp 1636968456
transform 1 0 46092 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_501
timestamp 1636968456
transform 1 0 47196 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_513
timestamp 1636968456
transform 1 0 48300 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_525
timestamp 1
transform 1 0 49404 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_531
timestamp 1
transform 1 0 49956 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_533
timestamp 1636968456
transform 1 0 50140 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_545
timestamp 1636968456
transform 1 0 51244 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_557
timestamp 1636968456
transform 1 0 52348 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_569
timestamp 1636968456
transform 1 0 53452 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_581
timestamp 1
transform 1 0 54556 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_587
timestamp 1
transform 1 0 55108 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_589
timestamp 1636968456
transform 1 0 55292 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_601
timestamp 1636968456
transform 1 0 56396 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_613
timestamp 1636968456
transform 1 0 57500 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_625
timestamp 1636968456
transform 1 0 58604 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_637
timestamp 1
transform 1 0 59708 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_643
timestamp 1
transform 1 0 60260 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_645
timestamp 1636968456
transform 1 0 60444 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_657
timestamp 1636968456
transform 1 0 61548 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_669
timestamp 1636968456
transform 1 0 62652 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_681
timestamp 1636968456
transform 1 0 63756 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_693
timestamp 1
transform 1 0 64860 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_699
timestamp 1
transform 1 0 65412 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_701
timestamp 1636968456
transform 1 0 65596 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_713
timestamp 1636968456
transform 1 0 66700 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_725
timestamp 1636968456
transform 1 0 67804 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_737
timestamp 1636968456
transform 1 0 68908 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_749
timestamp 1
transform 1 0 70012 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_755
timestamp 1
transform 1 0 70564 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_757
timestamp 1636968456
transform 1 0 70748 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_769
timestamp 1636968456
transform 1 0 71852 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_781
timestamp 1636968456
transform 1 0 72956 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_793
timestamp 1636968456
transform 1 0 74060 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_805
timestamp 1
transform 1 0 75164 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_811
timestamp 1
transform 1 0 75716 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_813
timestamp 1636968456
transform 1 0 75900 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_825
timestamp 1636968456
transform 1 0 77004 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_837
timestamp 1636968456
transform 1 0 78108 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_849
timestamp 1636968456
transform 1 0 79212 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_861
timestamp 1
transform 1 0 80316 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_867
timestamp 1
transform 1 0 80868 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_869
timestamp 1636968456
transform 1 0 81052 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_881
timestamp 1636968456
transform 1 0 82156 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_893
timestamp 1636968456
transform 1 0 83260 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_905
timestamp 1636968456
transform 1 0 84364 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_917
timestamp 1
transform 1 0 85468 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_923
timestamp 1
transform 1 0 86020 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_925
timestamp 1636968456
transform 1 0 86204 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_937
timestamp 1636968456
transform 1 0 87308 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_949
timestamp 1636968456
transform 1 0 88412 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_961
timestamp 1636968456
transform 1 0 89516 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_973
timestamp 1
transform 1 0 90620 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_979
timestamp 1
transform 1 0 91172 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_981
timestamp 1636968456
transform 1 0 91356 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_993
timestamp 1636968456
transform 1 0 92460 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_1005
timestamp 1636968456
transform 1 0 93564 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_1017
timestamp 1636968456
transform 1 0 94668 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_128_1029
timestamp 1
transform 1 0 95772 0 1 71808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_128_1035
timestamp 1
transform 1 0 96324 0 1 71808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_1037
timestamp 1636968456
transform 1 0 96508 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_1049
timestamp 1636968456
transform 1 0 97612 0 1 71808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_1061
timestamp 1636968456
transform 1 0 98716 0 1 71808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_128_1073
timestamp 1
transform 1 0 99820 0 1 71808
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_129_3
timestamp 1636968456
transform 1 0 1380 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_15
timestamp 1636968456
transform 1 0 2484 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_27
timestamp 1636968456
transform 1 0 3588 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_39
timestamp 1636968456
transform 1 0 4692 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_129_51
timestamp 1
transform 1 0 5796 0 -1 72896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_129_55
timestamp 1
transform 1 0 6164 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_57
timestamp 1636968456
transform 1 0 6348 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_69
timestamp 1636968456
transform 1 0 7452 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_81
timestamp 1636968456
transform 1 0 8556 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_93
timestamp 1636968456
transform 1 0 9660 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_105
timestamp 1
transform 1 0 10764 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_111
timestamp 1
transform 1 0 11316 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_113
timestamp 1636968456
transform 1 0 11500 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_125
timestamp 1636968456
transform 1 0 12604 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_137
timestamp 1636968456
transform 1 0 13708 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_149
timestamp 1636968456
transform 1 0 14812 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_161
timestamp 1
transform 1 0 15916 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_167
timestamp 1
transform 1 0 16468 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_169
timestamp 1636968456
transform 1 0 16652 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_181
timestamp 1636968456
transform 1 0 17756 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_193
timestamp 1636968456
transform 1 0 18860 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_205
timestamp 1636968456
transform 1 0 19964 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_217
timestamp 1
transform 1 0 21068 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_223
timestamp 1
transform 1 0 21620 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_225
timestamp 1636968456
transform 1 0 21804 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_237
timestamp 1636968456
transform 1 0 22908 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_249
timestamp 1636968456
transform 1 0 24012 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_261
timestamp 1636968456
transform 1 0 25116 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_273
timestamp 1
transform 1 0 26220 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_279
timestamp 1
transform 1 0 26772 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_281
timestamp 1636968456
transform 1 0 26956 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_293
timestamp 1636968456
transform 1 0 28060 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_305
timestamp 1636968456
transform 1 0 29164 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_317
timestamp 1636968456
transform 1 0 30268 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_329
timestamp 1
transform 1 0 31372 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_335
timestamp 1
transform 1 0 31924 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_337
timestamp 1636968456
transform 1 0 32108 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_349
timestamp 1636968456
transform 1 0 33212 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_361
timestamp 1636968456
transform 1 0 34316 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_373
timestamp 1636968456
transform 1 0 35420 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_385
timestamp 1
transform 1 0 36524 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_391
timestamp 1
transform 1 0 37076 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_393
timestamp 1636968456
transform 1 0 37260 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_405
timestamp 1636968456
transform 1 0 38364 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_417
timestamp 1636968456
transform 1 0 39468 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_429
timestamp 1636968456
transform 1 0 40572 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_441
timestamp 1
transform 1 0 41676 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_447
timestamp 1
transform 1 0 42228 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_449
timestamp 1636968456
transform 1 0 42412 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_461
timestamp 1636968456
transform 1 0 43516 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_473
timestamp 1636968456
transform 1 0 44620 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_485
timestamp 1636968456
transform 1 0 45724 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_497
timestamp 1
transform 1 0 46828 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_503
timestamp 1
transform 1 0 47380 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_505
timestamp 1636968456
transform 1 0 47564 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_517
timestamp 1636968456
transform 1 0 48668 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_529
timestamp 1636968456
transform 1 0 49772 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_541
timestamp 1636968456
transform 1 0 50876 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_553
timestamp 1
transform 1 0 51980 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_559
timestamp 1
transform 1 0 52532 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_561
timestamp 1636968456
transform 1 0 52716 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_573
timestamp 1636968456
transform 1 0 53820 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_585
timestamp 1636968456
transform 1 0 54924 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_597
timestamp 1636968456
transform 1 0 56028 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_609
timestamp 1
transform 1 0 57132 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_615
timestamp 1
transform 1 0 57684 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_617
timestamp 1636968456
transform 1 0 57868 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_629
timestamp 1636968456
transform 1 0 58972 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_641
timestamp 1636968456
transform 1 0 60076 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_653
timestamp 1636968456
transform 1 0 61180 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_665
timestamp 1
transform 1 0 62284 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_671
timestamp 1
transform 1 0 62836 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_673
timestamp 1636968456
transform 1 0 63020 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_685
timestamp 1636968456
transform 1 0 64124 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_697
timestamp 1636968456
transform 1 0 65228 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_709
timestamp 1636968456
transform 1 0 66332 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_721
timestamp 1
transform 1 0 67436 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_727
timestamp 1
transform 1 0 67988 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_729
timestamp 1636968456
transform 1 0 68172 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_741
timestamp 1636968456
transform 1 0 69276 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_753
timestamp 1636968456
transform 1 0 70380 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_765
timestamp 1636968456
transform 1 0 71484 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_777
timestamp 1
transform 1 0 72588 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_783
timestamp 1
transform 1 0 73140 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_785
timestamp 1636968456
transform 1 0 73324 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_797
timestamp 1636968456
transform 1 0 74428 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_809
timestamp 1636968456
transform 1 0 75532 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_821
timestamp 1636968456
transform 1 0 76636 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_833
timestamp 1
transform 1 0 77740 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_839
timestamp 1
transform 1 0 78292 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_841
timestamp 1636968456
transform 1 0 78476 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_853
timestamp 1636968456
transform 1 0 79580 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_865
timestamp 1636968456
transform 1 0 80684 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_877
timestamp 1636968456
transform 1 0 81788 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_889
timestamp 1
transform 1 0 82892 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_895
timestamp 1
transform 1 0 83444 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_897
timestamp 1636968456
transform 1 0 83628 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_909
timestamp 1636968456
transform 1 0 84732 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_921
timestamp 1636968456
transform 1 0 85836 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_933
timestamp 1636968456
transform 1 0 86940 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_945
timestamp 1
transform 1 0 88044 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_951
timestamp 1
transform 1 0 88596 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_953
timestamp 1636968456
transform 1 0 88780 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_965
timestamp 1636968456
transform 1 0 89884 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_977
timestamp 1636968456
transform 1 0 90988 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_989
timestamp 1636968456
transform 1 0 92092 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_1001
timestamp 1
transform 1 0 93196 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_1007
timestamp 1
transform 1 0 93748 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_1009
timestamp 1636968456
transform 1 0 93932 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_1021
timestamp 1636968456
transform 1 0 95036 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_1033
timestamp 1636968456
transform 1 0 96140 0 -1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_129_1045
timestamp 1636968456
transform 1 0 97244 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_129_1057
timestamp 1
transform 1 0 98348 0 -1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_129_1063
timestamp 1
transform 1 0 98900 0 -1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_1065
timestamp 1636968456
transform 1 0 99084 0 -1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_129_1077
timestamp 1
transform 1 0 100188 0 -1 72896
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_130_3
timestamp 1636968456
transform 1 0 1380 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_15
timestamp 1636968456
transform 1 0 2484 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_130_27
timestamp 1
transform 1 0 3588 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_29
timestamp 1636968456
transform 1 0 3772 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_41
timestamp 1636968456
transform 1 0 4876 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_53
timestamp 1636968456
transform 1 0 5980 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_65
timestamp 1636968456
transform 1 0 7084 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_77
timestamp 1
transform 1 0 8188 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_83
timestamp 1
transform 1 0 8740 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_85
timestamp 1636968456
transform 1 0 8924 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_97
timestamp 1636968456
transform 1 0 10028 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_109
timestamp 1636968456
transform 1 0 11132 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_121
timestamp 1636968456
transform 1 0 12236 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_133
timestamp 1
transform 1 0 13340 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_139
timestamp 1
transform 1 0 13892 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_141
timestamp 1636968456
transform 1 0 14076 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_153
timestamp 1636968456
transform 1 0 15180 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_165
timestamp 1636968456
transform 1 0 16284 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_177
timestamp 1636968456
transform 1 0 17388 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_189
timestamp 1
transform 1 0 18492 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_195
timestamp 1
transform 1 0 19044 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_197
timestamp 1636968456
transform 1 0 19228 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_209
timestamp 1636968456
transform 1 0 20332 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_221
timestamp 1636968456
transform 1 0 21436 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_233
timestamp 1636968456
transform 1 0 22540 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_245
timestamp 1
transform 1 0 23644 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_251
timestamp 1
transform 1 0 24196 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_253
timestamp 1636968456
transform 1 0 24380 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_265
timestamp 1636968456
transform 1 0 25484 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_277
timestamp 1636968456
transform 1 0 26588 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_289
timestamp 1636968456
transform 1 0 27692 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_301
timestamp 1
transform 1 0 28796 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_307
timestamp 1
transform 1 0 29348 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_309
timestamp 1636968456
transform 1 0 29532 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_321
timestamp 1636968456
transform 1 0 30636 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_333
timestamp 1636968456
transform 1 0 31740 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_345
timestamp 1636968456
transform 1 0 32844 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_357
timestamp 1
transform 1 0 33948 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_363
timestamp 1
transform 1 0 34500 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_365
timestamp 1636968456
transform 1 0 34684 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_377
timestamp 1636968456
transform 1 0 35788 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_389
timestamp 1636968456
transform 1 0 36892 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_401
timestamp 1636968456
transform 1 0 37996 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_413
timestamp 1
transform 1 0 39100 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_419
timestamp 1
transform 1 0 39652 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_421
timestamp 1636968456
transform 1 0 39836 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_433
timestamp 1636968456
transform 1 0 40940 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_445
timestamp 1636968456
transform 1 0 42044 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_457
timestamp 1636968456
transform 1 0 43148 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_469
timestamp 1
transform 1 0 44252 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_475
timestamp 1
transform 1 0 44804 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_477
timestamp 1636968456
transform 1 0 44988 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_489
timestamp 1636968456
transform 1 0 46092 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_501
timestamp 1636968456
transform 1 0 47196 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_513
timestamp 1636968456
transform 1 0 48300 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_525
timestamp 1
transform 1 0 49404 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_531
timestamp 1
transform 1 0 49956 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_533
timestamp 1636968456
transform 1 0 50140 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_545
timestamp 1636968456
transform 1 0 51244 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_557
timestamp 1636968456
transform 1 0 52348 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_569
timestamp 1636968456
transform 1 0 53452 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_581
timestamp 1
transform 1 0 54556 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_587
timestamp 1
transform 1 0 55108 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_589
timestamp 1636968456
transform 1 0 55292 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_601
timestamp 1636968456
transform 1 0 56396 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_613
timestamp 1636968456
transform 1 0 57500 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_625
timestamp 1636968456
transform 1 0 58604 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_637
timestamp 1
transform 1 0 59708 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_643
timestamp 1
transform 1 0 60260 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_645
timestamp 1636968456
transform 1 0 60444 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_657
timestamp 1636968456
transform 1 0 61548 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_669
timestamp 1636968456
transform 1 0 62652 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_681
timestamp 1636968456
transform 1 0 63756 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_693
timestamp 1
transform 1 0 64860 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_699
timestamp 1
transform 1 0 65412 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_701
timestamp 1636968456
transform 1 0 65596 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_713
timestamp 1636968456
transform 1 0 66700 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_725
timestamp 1636968456
transform 1 0 67804 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_737
timestamp 1636968456
transform 1 0 68908 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_749
timestamp 1
transform 1 0 70012 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_755
timestamp 1
transform 1 0 70564 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_757
timestamp 1636968456
transform 1 0 70748 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_769
timestamp 1636968456
transform 1 0 71852 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_781
timestamp 1636968456
transform 1 0 72956 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_793
timestamp 1636968456
transform 1 0 74060 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_805
timestamp 1
transform 1 0 75164 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_811
timestamp 1
transform 1 0 75716 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_813
timestamp 1636968456
transform 1 0 75900 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_825
timestamp 1636968456
transform 1 0 77004 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_837
timestamp 1636968456
transform 1 0 78108 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_849
timestamp 1636968456
transform 1 0 79212 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_861
timestamp 1
transform 1 0 80316 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_867
timestamp 1
transform 1 0 80868 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_869
timestamp 1636968456
transform 1 0 81052 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_881
timestamp 1636968456
transform 1 0 82156 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_893
timestamp 1636968456
transform 1 0 83260 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_905
timestamp 1636968456
transform 1 0 84364 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_917
timestamp 1
transform 1 0 85468 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_923
timestamp 1
transform 1 0 86020 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_925
timestamp 1636968456
transform 1 0 86204 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_937
timestamp 1636968456
transform 1 0 87308 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_949
timestamp 1636968456
transform 1 0 88412 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_961
timestamp 1636968456
transform 1 0 89516 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_973
timestamp 1
transform 1 0 90620 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_979
timestamp 1
transform 1 0 91172 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_981
timestamp 1636968456
transform 1 0 91356 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_993
timestamp 1636968456
transform 1 0 92460 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_1005
timestamp 1636968456
transform 1 0 93564 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_1017
timestamp 1636968456
transform 1 0 94668 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_130_1029
timestamp 1
transform 1 0 95772 0 1 72896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_130_1035
timestamp 1
transform 1 0 96324 0 1 72896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_1037
timestamp 1636968456
transform 1 0 96508 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_1049
timestamp 1636968456
transform 1 0 97612 0 1 72896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_130_1061
timestamp 1636968456
transform 1 0 98716 0 1 72896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_130_1073
timestamp 1
transform 1 0 99820 0 1 72896
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_131_3
timestamp 1636968456
transform 1 0 1380 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_15
timestamp 1636968456
transform 1 0 2484 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_27
timestamp 1636968456
transform 1 0 3588 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_39
timestamp 1636968456
transform 1 0 4692 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_131_51
timestamp 1
transform 1 0 5796 0 -1 73984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_131_55
timestamp 1
transform 1 0 6164 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_57
timestamp 1636968456
transform 1 0 6348 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_69
timestamp 1636968456
transform 1 0 7452 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_81
timestamp 1636968456
transform 1 0 8556 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_93
timestamp 1636968456
transform 1 0 9660 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_105
timestamp 1
transform 1 0 10764 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_111
timestamp 1
transform 1 0 11316 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_113
timestamp 1636968456
transform 1 0 11500 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_125
timestamp 1636968456
transform 1 0 12604 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_137
timestamp 1636968456
transform 1 0 13708 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_149
timestamp 1636968456
transform 1 0 14812 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_161
timestamp 1
transform 1 0 15916 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_167
timestamp 1
transform 1 0 16468 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_169
timestamp 1636968456
transform 1 0 16652 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_181
timestamp 1636968456
transform 1 0 17756 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_193
timestamp 1636968456
transform 1 0 18860 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_205
timestamp 1636968456
transform 1 0 19964 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_217
timestamp 1
transform 1 0 21068 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_223
timestamp 1
transform 1 0 21620 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_225
timestamp 1636968456
transform 1 0 21804 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_237
timestamp 1636968456
transform 1 0 22908 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_249
timestamp 1636968456
transform 1 0 24012 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_261
timestamp 1636968456
transform 1 0 25116 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_273
timestamp 1
transform 1 0 26220 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_279
timestamp 1
transform 1 0 26772 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_281
timestamp 1636968456
transform 1 0 26956 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_293
timestamp 1636968456
transform 1 0 28060 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_305
timestamp 1636968456
transform 1 0 29164 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_317
timestamp 1636968456
transform 1 0 30268 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_329
timestamp 1
transform 1 0 31372 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_335
timestamp 1
transform 1 0 31924 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_337
timestamp 1636968456
transform 1 0 32108 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_349
timestamp 1636968456
transform 1 0 33212 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_361
timestamp 1636968456
transform 1 0 34316 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_373
timestamp 1636968456
transform 1 0 35420 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_385
timestamp 1
transform 1 0 36524 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_391
timestamp 1
transform 1 0 37076 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_393
timestamp 1636968456
transform 1 0 37260 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_405
timestamp 1636968456
transform 1 0 38364 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_417
timestamp 1636968456
transform 1 0 39468 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_429
timestamp 1636968456
transform 1 0 40572 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_441
timestamp 1
transform 1 0 41676 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_447
timestamp 1
transform 1 0 42228 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_449
timestamp 1636968456
transform 1 0 42412 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_461
timestamp 1636968456
transform 1 0 43516 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_473
timestamp 1636968456
transform 1 0 44620 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_485
timestamp 1636968456
transform 1 0 45724 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_497
timestamp 1
transform 1 0 46828 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_503
timestamp 1
transform 1 0 47380 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_505
timestamp 1636968456
transform 1 0 47564 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_517
timestamp 1636968456
transform 1 0 48668 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_529
timestamp 1636968456
transform 1 0 49772 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_541
timestamp 1636968456
transform 1 0 50876 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_553
timestamp 1
transform 1 0 51980 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_559
timestamp 1
transform 1 0 52532 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_561
timestamp 1636968456
transform 1 0 52716 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_573
timestamp 1636968456
transform 1 0 53820 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_585
timestamp 1636968456
transform 1 0 54924 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_597
timestamp 1636968456
transform 1 0 56028 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_609
timestamp 1
transform 1 0 57132 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_615
timestamp 1
transform 1 0 57684 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_617
timestamp 1636968456
transform 1 0 57868 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_629
timestamp 1636968456
transform 1 0 58972 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_641
timestamp 1636968456
transform 1 0 60076 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_653
timestamp 1636968456
transform 1 0 61180 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_665
timestamp 1
transform 1 0 62284 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_671
timestamp 1
transform 1 0 62836 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_673
timestamp 1636968456
transform 1 0 63020 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_685
timestamp 1636968456
transform 1 0 64124 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_697
timestamp 1636968456
transform 1 0 65228 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_709
timestamp 1636968456
transform 1 0 66332 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_721
timestamp 1
transform 1 0 67436 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_727
timestamp 1
transform 1 0 67988 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_729
timestamp 1636968456
transform 1 0 68172 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_741
timestamp 1636968456
transform 1 0 69276 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_753
timestamp 1636968456
transform 1 0 70380 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_765
timestamp 1636968456
transform 1 0 71484 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_777
timestamp 1
transform 1 0 72588 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_783
timestamp 1
transform 1 0 73140 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_785
timestamp 1636968456
transform 1 0 73324 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_797
timestamp 1636968456
transform 1 0 74428 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_809
timestamp 1636968456
transform 1 0 75532 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_821
timestamp 1636968456
transform 1 0 76636 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_833
timestamp 1
transform 1 0 77740 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_839
timestamp 1
transform 1 0 78292 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_841
timestamp 1636968456
transform 1 0 78476 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_853
timestamp 1636968456
transform 1 0 79580 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_865
timestamp 1636968456
transform 1 0 80684 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_877
timestamp 1636968456
transform 1 0 81788 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_889
timestamp 1
transform 1 0 82892 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_895
timestamp 1
transform 1 0 83444 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_897
timestamp 1636968456
transform 1 0 83628 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_909
timestamp 1636968456
transform 1 0 84732 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_921
timestamp 1636968456
transform 1 0 85836 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_933
timestamp 1636968456
transform 1 0 86940 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_945
timestamp 1
transform 1 0 88044 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_951
timestamp 1
transform 1 0 88596 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_953
timestamp 1636968456
transform 1 0 88780 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_965
timestamp 1636968456
transform 1 0 89884 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_977
timestamp 1636968456
transform 1 0 90988 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_989
timestamp 1636968456
transform 1 0 92092 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_1001
timestamp 1
transform 1 0 93196 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_1007
timestamp 1
transform 1 0 93748 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_1009
timestamp 1636968456
transform 1 0 93932 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_1021
timestamp 1636968456
transform 1 0 95036 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_1033
timestamp 1636968456
transform 1 0 96140 0 -1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_1045
timestamp 1636968456
transform 1 0 97244 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_131_1057
timestamp 1
transform 1 0 98348 0 -1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_131_1063
timestamp 1
transform 1 0 98900 0 -1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_1065
timestamp 1636968456
transform 1 0 99084 0 -1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_131_1077
timestamp 1
transform 1 0 100188 0 -1 73984
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_132_3
timestamp 1636968456
transform 1 0 1380 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_15
timestamp 1636968456
transform 1 0 2484 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_132_27
timestamp 1
transform 1 0 3588 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_29
timestamp 1636968456
transform 1 0 3772 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_41
timestamp 1636968456
transform 1 0 4876 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_53
timestamp 1636968456
transform 1 0 5980 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_65
timestamp 1636968456
transform 1 0 7084 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_77
timestamp 1
transform 1 0 8188 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_83
timestamp 1
transform 1 0 8740 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_85
timestamp 1636968456
transform 1 0 8924 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_97
timestamp 1636968456
transform 1 0 10028 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_109
timestamp 1636968456
transform 1 0 11132 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_121
timestamp 1636968456
transform 1 0 12236 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_133
timestamp 1
transform 1 0 13340 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_139
timestamp 1
transform 1 0 13892 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_141
timestamp 1636968456
transform 1 0 14076 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_153
timestamp 1636968456
transform 1 0 15180 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_165
timestamp 1636968456
transform 1 0 16284 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_177
timestamp 1636968456
transform 1 0 17388 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_189
timestamp 1
transform 1 0 18492 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_195
timestamp 1
transform 1 0 19044 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_197
timestamp 1636968456
transform 1 0 19228 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_209
timestamp 1636968456
transform 1 0 20332 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_221
timestamp 1636968456
transform 1 0 21436 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_233
timestamp 1636968456
transform 1 0 22540 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_245
timestamp 1
transform 1 0 23644 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_251
timestamp 1
transform 1 0 24196 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_253
timestamp 1636968456
transform 1 0 24380 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_265
timestamp 1636968456
transform 1 0 25484 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_277
timestamp 1636968456
transform 1 0 26588 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_289
timestamp 1636968456
transform 1 0 27692 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_301
timestamp 1
transform 1 0 28796 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_307
timestamp 1
transform 1 0 29348 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_309
timestamp 1636968456
transform 1 0 29532 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_321
timestamp 1636968456
transform 1 0 30636 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_333
timestamp 1636968456
transform 1 0 31740 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_345
timestamp 1636968456
transform 1 0 32844 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_357
timestamp 1
transform 1 0 33948 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_363
timestamp 1
transform 1 0 34500 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_365
timestamp 1636968456
transform 1 0 34684 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_377
timestamp 1636968456
transform 1 0 35788 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_389
timestamp 1636968456
transform 1 0 36892 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_401
timestamp 1636968456
transform 1 0 37996 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_413
timestamp 1
transform 1 0 39100 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_419
timestamp 1
transform 1 0 39652 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_421
timestamp 1636968456
transform 1 0 39836 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_433
timestamp 1636968456
transform 1 0 40940 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_445
timestamp 1636968456
transform 1 0 42044 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_457
timestamp 1636968456
transform 1 0 43148 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_469
timestamp 1
transform 1 0 44252 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_475
timestamp 1
transform 1 0 44804 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_477
timestamp 1636968456
transform 1 0 44988 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_489
timestamp 1636968456
transform 1 0 46092 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_501
timestamp 1636968456
transform 1 0 47196 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_513
timestamp 1636968456
transform 1 0 48300 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_525
timestamp 1
transform 1 0 49404 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_531
timestamp 1
transform 1 0 49956 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_533
timestamp 1636968456
transform 1 0 50140 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_545
timestamp 1636968456
transform 1 0 51244 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_557
timestamp 1636968456
transform 1 0 52348 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_569
timestamp 1636968456
transform 1 0 53452 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_581
timestamp 1
transform 1 0 54556 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_587
timestamp 1
transform 1 0 55108 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_589
timestamp 1636968456
transform 1 0 55292 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_601
timestamp 1636968456
transform 1 0 56396 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_613
timestamp 1636968456
transform 1 0 57500 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_625
timestamp 1636968456
transform 1 0 58604 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_637
timestamp 1
transform 1 0 59708 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_643
timestamp 1
transform 1 0 60260 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_645
timestamp 1636968456
transform 1 0 60444 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_657
timestamp 1636968456
transform 1 0 61548 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_669
timestamp 1636968456
transform 1 0 62652 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_681
timestamp 1636968456
transform 1 0 63756 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_693
timestamp 1
transform 1 0 64860 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_699
timestamp 1
transform 1 0 65412 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_701
timestamp 1636968456
transform 1 0 65596 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_713
timestamp 1636968456
transform 1 0 66700 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_725
timestamp 1636968456
transform 1 0 67804 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_737
timestamp 1636968456
transform 1 0 68908 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_749
timestamp 1
transform 1 0 70012 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_755
timestamp 1
transform 1 0 70564 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_757
timestamp 1636968456
transform 1 0 70748 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_769
timestamp 1636968456
transform 1 0 71852 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_781
timestamp 1636968456
transform 1 0 72956 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_793
timestamp 1636968456
transform 1 0 74060 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_805
timestamp 1
transform 1 0 75164 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_811
timestamp 1
transform 1 0 75716 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_813
timestamp 1636968456
transform 1 0 75900 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_825
timestamp 1636968456
transform 1 0 77004 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_837
timestamp 1636968456
transform 1 0 78108 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_849
timestamp 1636968456
transform 1 0 79212 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_861
timestamp 1
transform 1 0 80316 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_867
timestamp 1
transform 1 0 80868 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_869
timestamp 1636968456
transform 1 0 81052 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_881
timestamp 1636968456
transform 1 0 82156 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_893
timestamp 1636968456
transform 1 0 83260 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_905
timestamp 1636968456
transform 1 0 84364 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_917
timestamp 1
transform 1 0 85468 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_923
timestamp 1
transform 1 0 86020 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_925
timestamp 1636968456
transform 1 0 86204 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_937
timestamp 1636968456
transform 1 0 87308 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_949
timestamp 1636968456
transform 1 0 88412 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_961
timestamp 1636968456
transform 1 0 89516 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_973
timestamp 1
transform 1 0 90620 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_979
timestamp 1
transform 1 0 91172 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_981
timestamp 1636968456
transform 1 0 91356 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_993
timestamp 1636968456
transform 1 0 92460 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_1005
timestamp 1636968456
transform 1 0 93564 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_1017
timestamp 1636968456
transform 1 0 94668 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_132_1029
timestamp 1
transform 1 0 95772 0 1 73984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_132_1035
timestamp 1
transform 1 0 96324 0 1 73984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_1037
timestamp 1636968456
transform 1 0 96508 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_1049
timestamp 1636968456
transform 1 0 97612 0 1 73984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_1061
timestamp 1636968456
transform 1 0 98716 0 1 73984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_132_1073
timestamp 1
transform 1 0 99820 0 1 73984
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_133_3
timestamp 1636968456
transform 1 0 1380 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_15
timestamp 1636968456
transform 1 0 2484 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_27
timestamp 1636968456
transform 1 0 3588 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_39
timestamp 1636968456
transform 1 0 4692 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_133_51
timestamp 1
transform 1 0 5796 0 -1 75072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_133_55
timestamp 1
transform 1 0 6164 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_57
timestamp 1636968456
transform 1 0 6348 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_69
timestamp 1636968456
transform 1 0 7452 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_81
timestamp 1636968456
transform 1 0 8556 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_93
timestamp 1636968456
transform 1 0 9660 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_105
timestamp 1
transform 1 0 10764 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_111
timestamp 1
transform 1 0 11316 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_113
timestamp 1636968456
transform 1 0 11500 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_125
timestamp 1636968456
transform 1 0 12604 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_137
timestamp 1636968456
transform 1 0 13708 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_149
timestamp 1636968456
transform 1 0 14812 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_161
timestamp 1
transform 1 0 15916 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_167
timestamp 1
transform 1 0 16468 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_169
timestamp 1636968456
transform 1 0 16652 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_181
timestamp 1636968456
transform 1 0 17756 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_193
timestamp 1636968456
transform 1 0 18860 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_205
timestamp 1636968456
transform 1 0 19964 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_217
timestamp 1
transform 1 0 21068 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_223
timestamp 1
transform 1 0 21620 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_225
timestamp 1636968456
transform 1 0 21804 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_237
timestamp 1636968456
transform 1 0 22908 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_249
timestamp 1636968456
transform 1 0 24012 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_261
timestamp 1636968456
transform 1 0 25116 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_273
timestamp 1
transform 1 0 26220 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_279
timestamp 1
transform 1 0 26772 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_281
timestamp 1636968456
transform 1 0 26956 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_293
timestamp 1636968456
transform 1 0 28060 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_305
timestamp 1636968456
transform 1 0 29164 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_317
timestamp 1636968456
transform 1 0 30268 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_329
timestamp 1
transform 1 0 31372 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_335
timestamp 1
transform 1 0 31924 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_337
timestamp 1636968456
transform 1 0 32108 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_349
timestamp 1636968456
transform 1 0 33212 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_361
timestamp 1636968456
transform 1 0 34316 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_373
timestamp 1636968456
transform 1 0 35420 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_385
timestamp 1
transform 1 0 36524 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_391
timestamp 1
transform 1 0 37076 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_393
timestamp 1636968456
transform 1 0 37260 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_405
timestamp 1636968456
transform 1 0 38364 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_417
timestamp 1636968456
transform 1 0 39468 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_429
timestamp 1636968456
transform 1 0 40572 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_441
timestamp 1
transform 1 0 41676 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_447
timestamp 1
transform 1 0 42228 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_449
timestamp 1636968456
transform 1 0 42412 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_461
timestamp 1636968456
transform 1 0 43516 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_473
timestamp 1636968456
transform 1 0 44620 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_133_485
timestamp 1
transform 1 0 45724 0 -1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_133_496
timestamp 1
transform 1 0 46736 0 -1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_133_505
timestamp 1
transform 1 0 47564 0 -1 75072
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_133_514
timestamp 1636968456
transform 1 0 48392 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_133_526
timestamp 1
transform 1 0 49496 0 -1 75072
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_133_533
timestamp 1636968456
transform 1 0 50140 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_545
timestamp 1
transform 1 0 51244 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_133_554
timestamp 1
transform 1 0 52072 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_133_561
timestamp 1
transform 1 0 52716 0 -1 75072
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_133_568
timestamp 1636968456
transform 1 0 53360 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_133_580
timestamp 1
transform 1 0 54464 0 -1 75072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_133_586
timestamp 1636968456
transform 1 0 55016 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_598
timestamp 1
transform 1 0 56120 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_604
timestamp 1
transform 1 0 56672 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_133_608
timestamp 1
transform 1 0 57040 0 -1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_133_617
timestamp 1
transform 1 0 57868 0 -1 75072
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_133_624
timestamp 1636968456
transform 1 0 58512 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_133_636
timestamp 1
transform 1 0 59616 0 -1 75072
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_133_649
timestamp 1636968456
transform 1 0 60812 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_133_661
timestamp 1
transform 1 0 61916 0 -1 75072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_133_669
timestamp 1
transform 1 0 62652 0 -1 75072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_133_673
timestamp 1636968456
transform 1 0 63020 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_685
timestamp 1636968456
transform 1 0 64124 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_697
timestamp 1636968456
transform 1 0 65228 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_709
timestamp 1636968456
transform 1 0 66332 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_721
timestamp 1
transform 1 0 67436 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_727
timestamp 1
transform 1 0 67988 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_729
timestamp 1636968456
transform 1 0 68172 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_741
timestamp 1636968456
transform 1 0 69276 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_753
timestamp 1636968456
transform 1 0 70380 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_765
timestamp 1636968456
transform 1 0 71484 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_777
timestamp 1
transform 1 0 72588 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_783
timestamp 1
transform 1 0 73140 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_785
timestamp 1636968456
transform 1 0 73324 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_797
timestamp 1636968456
transform 1 0 74428 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_809
timestamp 1636968456
transform 1 0 75532 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_821
timestamp 1636968456
transform 1 0 76636 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_833
timestamp 1
transform 1 0 77740 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_839
timestamp 1
transform 1 0 78292 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_841
timestamp 1636968456
transform 1 0 78476 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_853
timestamp 1636968456
transform 1 0 79580 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_865
timestamp 1636968456
transform 1 0 80684 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_877
timestamp 1636968456
transform 1 0 81788 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_889
timestamp 1
transform 1 0 82892 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_895
timestamp 1
transform 1 0 83444 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_897
timestamp 1636968456
transform 1 0 83628 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_909
timestamp 1636968456
transform 1 0 84732 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_921
timestamp 1636968456
transform 1 0 85836 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_933
timestamp 1636968456
transform 1 0 86940 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_945
timestamp 1
transform 1 0 88044 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_951
timestamp 1
transform 1 0 88596 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_953
timestamp 1636968456
transform 1 0 88780 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_965
timestamp 1636968456
transform 1 0 89884 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_977
timestamp 1636968456
transform 1 0 90988 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_989
timestamp 1636968456
transform 1 0 92092 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_1001
timestamp 1
transform 1 0 93196 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_1007
timestamp 1
transform 1 0 93748 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_1009
timestamp 1636968456
transform 1 0 93932 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_1021
timestamp 1636968456
transform 1 0 95036 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_1033
timestamp 1636968456
transform 1 0 96140 0 -1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_133_1045
timestamp 1636968456
transform 1 0 97244 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_133_1057
timestamp 1
transform 1 0 98348 0 -1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_133_1063
timestamp 1
transform 1 0 98900 0 -1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_1065
timestamp 1636968456
transform 1 0 99084 0 -1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_133_1077
timestamp 1
transform 1 0 100188 0 -1 75072
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_134_3
timestamp 1636968456
transform 1 0 1380 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_15
timestamp 1636968456
transform 1 0 2484 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_134_27
timestamp 1
transform 1 0 3588 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_29
timestamp 1636968456
transform 1 0 3772 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_41
timestamp 1636968456
transform 1 0 4876 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_53
timestamp 1636968456
transform 1 0 5980 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_65
timestamp 1636968456
transform 1 0 7084 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_77
timestamp 1
transform 1 0 8188 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_83
timestamp 1
transform 1 0 8740 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_85
timestamp 1636968456
transform 1 0 8924 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_97
timestamp 1636968456
transform 1 0 10028 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_109
timestamp 1636968456
transform 1 0 11132 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_121
timestamp 1636968456
transform 1 0 12236 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_133
timestamp 1
transform 1 0 13340 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_139
timestamp 1
transform 1 0 13892 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_141
timestamp 1636968456
transform 1 0 14076 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_153
timestamp 1636968456
transform 1 0 15180 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_165
timestamp 1636968456
transform 1 0 16284 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_177
timestamp 1636968456
transform 1 0 17388 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_189
timestamp 1
transform 1 0 18492 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_195
timestamp 1
transform 1 0 19044 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_197
timestamp 1636968456
transform 1 0 19228 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_209
timestamp 1636968456
transform 1 0 20332 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_221
timestamp 1636968456
transform 1 0 21436 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_233
timestamp 1636968456
transform 1 0 22540 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_245
timestamp 1
transform 1 0 23644 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_251
timestamp 1
transform 1 0 24196 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_253
timestamp 1636968456
transform 1 0 24380 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_265
timestamp 1636968456
transform 1 0 25484 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_277
timestamp 1636968456
transform 1 0 26588 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_289
timestamp 1636968456
transform 1 0 27692 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_301
timestamp 1
transform 1 0 28796 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_307
timestamp 1
transform 1 0 29348 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_309
timestamp 1636968456
transform 1 0 29532 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_321
timestamp 1636968456
transform 1 0 30636 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_333
timestamp 1636968456
transform 1 0 31740 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_345
timestamp 1636968456
transform 1 0 32844 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_357
timestamp 1
transform 1 0 33948 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_363
timestamp 1
transform 1 0 34500 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_365
timestamp 1636968456
transform 1 0 34684 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_377
timestamp 1636968456
transform 1 0 35788 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_389
timestamp 1636968456
transform 1 0 36892 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_401
timestamp 1636968456
transform 1 0 37996 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_413
timestamp 1
transform 1 0 39100 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_419
timestamp 1
transform 1 0 39652 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_421
timestamp 1636968456
transform 1 0 39836 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_433
timestamp 1636968456
transform 1 0 40940 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_445
timestamp 1636968456
transform 1 0 42044 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_457
timestamp 1636968456
transform 1 0 43148 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_469
timestamp 1
transform 1 0 44252 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_475
timestamp 1
transform 1 0 44804 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_477
timestamp 1636968456
transform 1 0 44988 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_489
timestamp 1636968456
transform 1 0 46092 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_501
timestamp 1636968456
transform 1 0 47196 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_513
timestamp 1636968456
transform 1 0 48300 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_525
timestamp 1
transform 1 0 49404 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_531
timestamp 1
transform 1 0 49956 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_533
timestamp 1636968456
transform 1 0 50140 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_545
timestamp 1636968456
transform 1 0 51244 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_557
timestamp 1636968456
transform 1 0 52348 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_569
timestamp 1636968456
transform 1 0 53452 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_581
timestamp 1
transform 1 0 54556 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_587
timestamp 1
transform 1 0 55108 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_589
timestamp 1636968456
transform 1 0 55292 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_601
timestamp 1636968456
transform 1 0 56396 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_613
timestamp 1636968456
transform 1 0 57500 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_625
timestamp 1636968456
transform 1 0 58604 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_637
timestamp 1
transform 1 0 59708 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_643
timestamp 1
transform 1 0 60260 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_645
timestamp 1636968456
transform 1 0 60444 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_657
timestamp 1636968456
transform 1 0 61548 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_669
timestamp 1636968456
transform 1 0 62652 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_681
timestamp 1636968456
transform 1 0 63756 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_693
timestamp 1
transform 1 0 64860 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_699
timestamp 1
transform 1 0 65412 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_701
timestamp 1636968456
transform 1 0 65596 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_713
timestamp 1636968456
transform 1 0 66700 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_725
timestamp 1636968456
transform 1 0 67804 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_737
timestamp 1636968456
transform 1 0 68908 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_749
timestamp 1
transform 1 0 70012 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_755
timestamp 1
transform 1 0 70564 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_757
timestamp 1636968456
transform 1 0 70748 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_769
timestamp 1636968456
transform 1 0 71852 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_781
timestamp 1636968456
transform 1 0 72956 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_793
timestamp 1636968456
transform 1 0 74060 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_805
timestamp 1
transform 1 0 75164 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_811
timestamp 1
transform 1 0 75716 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_813
timestamp 1636968456
transform 1 0 75900 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_825
timestamp 1636968456
transform 1 0 77004 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_837
timestamp 1636968456
transform 1 0 78108 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_849
timestamp 1636968456
transform 1 0 79212 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_861
timestamp 1
transform 1 0 80316 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_867
timestamp 1
transform 1 0 80868 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_869
timestamp 1636968456
transform 1 0 81052 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_881
timestamp 1636968456
transform 1 0 82156 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_893
timestamp 1636968456
transform 1 0 83260 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_905
timestamp 1636968456
transform 1 0 84364 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_917
timestamp 1
transform 1 0 85468 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_923
timestamp 1
transform 1 0 86020 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_925
timestamp 1636968456
transform 1 0 86204 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_937
timestamp 1636968456
transform 1 0 87308 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_949
timestamp 1636968456
transform 1 0 88412 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_961
timestamp 1636968456
transform 1 0 89516 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_973
timestamp 1
transform 1 0 90620 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_979
timestamp 1
transform 1 0 91172 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_981
timestamp 1636968456
transform 1 0 91356 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_993
timestamp 1636968456
transform 1 0 92460 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_1005
timestamp 1636968456
transform 1 0 93564 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_1017
timestamp 1636968456
transform 1 0 94668 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_134_1029
timestamp 1
transform 1 0 95772 0 1 75072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_1035
timestamp 1
transform 1 0 96324 0 1 75072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_1037
timestamp 1636968456
transform 1 0 96508 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_1049
timestamp 1636968456
transform 1 0 97612 0 1 75072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_1061
timestamp 1636968456
transform 1 0 98716 0 1 75072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_134_1073
timestamp 1
transform 1 0 99820 0 1 75072
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_135_3
timestamp 1636968456
transform 1 0 1380 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_15
timestamp 1636968456
transform 1 0 2484 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_27
timestamp 1636968456
transform 1 0 3588 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_39
timestamp 1636968456
transform 1 0 4692 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_135_51
timestamp 1
transform 1 0 5796 0 -1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_135_55
timestamp 1
transform 1 0 6164 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_57
timestamp 1636968456
transform 1 0 6348 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_69
timestamp 1636968456
transform 1 0 7452 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_81
timestamp 1636968456
transform 1 0 8556 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_93
timestamp 1636968456
transform 1 0 9660 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_105
timestamp 1
transform 1 0 10764 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_111
timestamp 1
transform 1 0 11316 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_113
timestamp 1636968456
transform 1 0 11500 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_125
timestamp 1636968456
transform 1 0 12604 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_137
timestamp 1636968456
transform 1 0 13708 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_149
timestamp 1636968456
transform 1 0 14812 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_161
timestamp 1
transform 1 0 15916 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_167
timestamp 1
transform 1 0 16468 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_169
timestamp 1636968456
transform 1 0 16652 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_181
timestamp 1636968456
transform 1 0 17756 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_193
timestamp 1636968456
transform 1 0 18860 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_205
timestamp 1636968456
transform 1 0 19964 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_217
timestamp 1
transform 1 0 21068 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_223
timestamp 1
transform 1 0 21620 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_225
timestamp 1636968456
transform 1 0 21804 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_237
timestamp 1636968456
transform 1 0 22908 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_249
timestamp 1636968456
transform 1 0 24012 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_261
timestamp 1636968456
transform 1 0 25116 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_273
timestamp 1
transform 1 0 26220 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_279
timestamp 1
transform 1 0 26772 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_281
timestamp 1636968456
transform 1 0 26956 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_293
timestamp 1636968456
transform 1 0 28060 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_305
timestamp 1636968456
transform 1 0 29164 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_317
timestamp 1636968456
transform 1 0 30268 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_329
timestamp 1
transform 1 0 31372 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_335
timestamp 1
transform 1 0 31924 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_337
timestamp 1636968456
transform 1 0 32108 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_349
timestamp 1636968456
transform 1 0 33212 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_361
timestamp 1636968456
transform 1 0 34316 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_373
timestamp 1636968456
transform 1 0 35420 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_385
timestamp 1
transform 1 0 36524 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_391
timestamp 1
transform 1 0 37076 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_393
timestamp 1636968456
transform 1 0 37260 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_405
timestamp 1636968456
transform 1 0 38364 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_417
timestamp 1636968456
transform 1 0 39468 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_429
timestamp 1636968456
transform 1 0 40572 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_441
timestamp 1
transform 1 0 41676 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_447
timestamp 1
transform 1 0 42228 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_449
timestamp 1636968456
transform 1 0 42412 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_461
timestamp 1636968456
transform 1 0 43516 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_473
timestamp 1636968456
transform 1 0 44620 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_485
timestamp 1636968456
transform 1 0 45724 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_497
timestamp 1
transform 1 0 46828 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_503
timestamp 1
transform 1 0 47380 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_505
timestamp 1636968456
transform 1 0 47564 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_517
timestamp 1636968456
transform 1 0 48668 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_529
timestamp 1636968456
transform 1 0 49772 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_541
timestamp 1636968456
transform 1 0 50876 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_553
timestamp 1
transform 1 0 51980 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_559
timestamp 1
transform 1 0 52532 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_561
timestamp 1636968456
transform 1 0 52716 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_573
timestamp 1636968456
transform 1 0 53820 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_585
timestamp 1636968456
transform 1 0 54924 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_597
timestamp 1636968456
transform 1 0 56028 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_609
timestamp 1
transform 1 0 57132 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_615
timestamp 1
transform 1 0 57684 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_617
timestamp 1636968456
transform 1 0 57868 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_629
timestamp 1636968456
transform 1 0 58972 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_641
timestamp 1636968456
transform 1 0 60076 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_653
timestamp 1636968456
transform 1 0 61180 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_665
timestamp 1
transform 1 0 62284 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_671
timestamp 1
transform 1 0 62836 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_673
timestamp 1636968456
transform 1 0 63020 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_685
timestamp 1636968456
transform 1 0 64124 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_697
timestamp 1636968456
transform 1 0 65228 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_709
timestamp 1636968456
transform 1 0 66332 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_721
timestamp 1
transform 1 0 67436 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_727
timestamp 1
transform 1 0 67988 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_729
timestamp 1636968456
transform 1 0 68172 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_741
timestamp 1636968456
transform 1 0 69276 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_753
timestamp 1636968456
transform 1 0 70380 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_765
timestamp 1636968456
transform 1 0 71484 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_777
timestamp 1
transform 1 0 72588 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_783
timestamp 1
transform 1 0 73140 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_785
timestamp 1636968456
transform 1 0 73324 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_797
timestamp 1636968456
transform 1 0 74428 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_809
timestamp 1636968456
transform 1 0 75532 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_821
timestamp 1636968456
transform 1 0 76636 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_833
timestamp 1
transform 1 0 77740 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_839
timestamp 1
transform 1 0 78292 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_841
timestamp 1636968456
transform 1 0 78476 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_853
timestamp 1636968456
transform 1 0 79580 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_865
timestamp 1636968456
transform 1 0 80684 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_877
timestamp 1636968456
transform 1 0 81788 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_889
timestamp 1
transform 1 0 82892 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_895
timestamp 1
transform 1 0 83444 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_897
timestamp 1636968456
transform 1 0 83628 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_909
timestamp 1636968456
transform 1 0 84732 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_921
timestamp 1636968456
transform 1 0 85836 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_933
timestamp 1636968456
transform 1 0 86940 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_945
timestamp 1
transform 1 0 88044 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_951
timestamp 1
transform 1 0 88596 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_953
timestamp 1636968456
transform 1 0 88780 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_965
timestamp 1636968456
transform 1 0 89884 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_977
timestamp 1636968456
transform 1 0 90988 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_989
timestamp 1636968456
transform 1 0 92092 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_1001
timestamp 1
transform 1 0 93196 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_1007
timestamp 1
transform 1 0 93748 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_1009
timestamp 1636968456
transform 1 0 93932 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_1021
timestamp 1636968456
transform 1 0 95036 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_1033
timestamp 1636968456
transform 1 0 96140 0 -1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_135_1045
timestamp 1636968456
transform 1 0 97244 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_135_1057
timestamp 1
transform 1 0 98348 0 -1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_135_1063
timestamp 1
transform 1 0 98900 0 -1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_1065
timestamp 1636968456
transform 1 0 99084 0 -1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_135_1077
timestamp 1
transform 1 0 100188 0 -1 76160
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_136_3
timestamp 1636968456
transform 1 0 1380 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_15
timestamp 1636968456
transform 1 0 2484 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_136_27
timestamp 1
transform 1 0 3588 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_29
timestamp 1636968456
transform 1 0 3772 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_41
timestamp 1636968456
transform 1 0 4876 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_53
timestamp 1636968456
transform 1 0 5980 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_65
timestamp 1636968456
transform 1 0 7084 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_77
timestamp 1
transform 1 0 8188 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_83
timestamp 1
transform 1 0 8740 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_85
timestamp 1636968456
transform 1 0 8924 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_97
timestamp 1636968456
transform 1 0 10028 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_109
timestamp 1636968456
transform 1 0 11132 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_121
timestamp 1636968456
transform 1 0 12236 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_133
timestamp 1
transform 1 0 13340 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_139
timestamp 1
transform 1 0 13892 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_141
timestamp 1636968456
transform 1 0 14076 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_153
timestamp 1636968456
transform 1 0 15180 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_165
timestamp 1636968456
transform 1 0 16284 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_177
timestamp 1636968456
transform 1 0 17388 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_189
timestamp 1
transform 1 0 18492 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_195
timestamp 1
transform 1 0 19044 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_197
timestamp 1636968456
transform 1 0 19228 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_209
timestamp 1636968456
transform 1 0 20332 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_221
timestamp 1636968456
transform 1 0 21436 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_233
timestamp 1636968456
transform 1 0 22540 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_245
timestamp 1
transform 1 0 23644 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_251
timestamp 1
transform 1 0 24196 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_253
timestamp 1636968456
transform 1 0 24380 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_265
timestamp 1636968456
transform 1 0 25484 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_277
timestamp 1636968456
transform 1 0 26588 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_289
timestamp 1636968456
transform 1 0 27692 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_301
timestamp 1
transform 1 0 28796 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_307
timestamp 1
transform 1 0 29348 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_309
timestamp 1636968456
transform 1 0 29532 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_321
timestamp 1636968456
transform 1 0 30636 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_333
timestamp 1636968456
transform 1 0 31740 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_345
timestamp 1636968456
transform 1 0 32844 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_357
timestamp 1
transform 1 0 33948 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_363
timestamp 1
transform 1 0 34500 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_365
timestamp 1636968456
transform 1 0 34684 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_377
timestamp 1636968456
transform 1 0 35788 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_389
timestamp 1636968456
transform 1 0 36892 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_401
timestamp 1636968456
transform 1 0 37996 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_413
timestamp 1
transform 1 0 39100 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_419
timestamp 1
transform 1 0 39652 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_421
timestamp 1636968456
transform 1 0 39836 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_433
timestamp 1636968456
transform 1 0 40940 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_445
timestamp 1636968456
transform 1 0 42044 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_136_457
timestamp 1
transform 1 0 43148 0 1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_136_461
timestamp 1
transform 1 0 43516 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_464
timestamp 1636968456
transform 1 0 43792 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_477
timestamp 1636968456
transform 1 0 44988 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_489
timestamp 1636968456
transform 1 0 46092 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_501
timestamp 1636968456
transform 1 0 47196 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_513
timestamp 1636968456
transform 1 0 48300 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_136_527
timestamp 1
transform 1 0 49588 0 1 76160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_136_531
timestamp 1
transform 1 0 49956 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_533
timestamp 1636968456
transform 1 0 50140 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_545
timestamp 1636968456
transform 1 0 51244 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_557
timestamp 1636968456
transform 1 0 52348 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_569
timestamp 1636968456
transform 1 0 53452 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_581
timestamp 1
transform 1 0 54556 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_587
timestamp 1
transform 1 0 55108 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_589
timestamp 1636968456
transform 1 0 55292 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_601
timestamp 1636968456
transform 1 0 56396 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_613
timestamp 1636968456
transform 1 0 57500 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_625
timestamp 1636968456
transform 1 0 58604 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_637
timestamp 1
transform 1 0 59708 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_643
timestamp 1
transform 1 0 60260 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_645
timestamp 1636968456
transform 1 0 60444 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_657
timestamp 1636968456
transform 1 0 61548 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_669
timestamp 1636968456
transform 1 0 62652 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_681
timestamp 1636968456
transform 1 0 63756 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_693
timestamp 1
transform 1 0 64860 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_699
timestamp 1
transform 1 0 65412 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_701
timestamp 1636968456
transform 1 0 65596 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_713
timestamp 1636968456
transform 1 0 66700 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_725
timestamp 1636968456
transform 1 0 67804 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_737
timestamp 1636968456
transform 1 0 68908 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_749
timestamp 1
transform 1 0 70012 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_755
timestamp 1
transform 1 0 70564 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_757
timestamp 1636968456
transform 1 0 70748 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_769
timestamp 1636968456
transform 1 0 71852 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_781
timestamp 1636968456
transform 1 0 72956 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_793
timestamp 1636968456
transform 1 0 74060 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_805
timestamp 1
transform 1 0 75164 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_811
timestamp 1
transform 1 0 75716 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_813
timestamp 1636968456
transform 1 0 75900 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_825
timestamp 1636968456
transform 1 0 77004 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_837
timestamp 1636968456
transform 1 0 78108 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_849
timestamp 1636968456
transform 1 0 79212 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_861
timestamp 1
transform 1 0 80316 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_867
timestamp 1
transform 1 0 80868 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_869
timestamp 1636968456
transform 1 0 81052 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_881
timestamp 1636968456
transform 1 0 82156 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_893
timestamp 1636968456
transform 1 0 83260 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_905
timestamp 1636968456
transform 1 0 84364 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_917
timestamp 1
transform 1 0 85468 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_923
timestamp 1
transform 1 0 86020 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_925
timestamp 1636968456
transform 1 0 86204 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_937
timestamp 1636968456
transform 1 0 87308 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_949
timestamp 1636968456
transform 1 0 88412 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_961
timestamp 1636968456
transform 1 0 89516 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_973
timestamp 1
transform 1 0 90620 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_979
timestamp 1
transform 1 0 91172 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_981
timestamp 1636968456
transform 1 0 91356 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_993
timestamp 1636968456
transform 1 0 92460 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_1005
timestamp 1636968456
transform 1 0 93564 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_1017
timestamp 1636968456
transform 1 0 94668 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_1029
timestamp 1
transform 1 0 95772 0 1 76160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_136_1035
timestamp 1
transform 1 0 96324 0 1 76160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_1037
timestamp 1636968456
transform 1 0 96508 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_1049
timestamp 1636968456
transform 1 0 97612 0 1 76160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_1061
timestamp 1636968456
transform 1 0 98716 0 1 76160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_136_1073
timestamp 1
transform 1 0 99820 0 1 76160
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_137_3
timestamp 1636968456
transform 1 0 1380 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_15
timestamp 1636968456
transform 1 0 2484 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_27
timestamp 1636968456
transform 1 0 3588 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_39
timestamp 1636968456
transform 1 0 4692 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_137_51
timestamp 1
transform 1 0 5796 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_137_55
timestamp 1
transform 1 0 6164 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_57
timestamp 1636968456
transform 1 0 6348 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_69
timestamp 1636968456
transform 1 0 7452 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_81
timestamp 1636968456
transform 1 0 8556 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_93
timestamp 1636968456
transform 1 0 9660 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_105
timestamp 1
transform 1 0 10764 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_111
timestamp 1
transform 1 0 11316 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_113
timestamp 1636968456
transform 1 0 11500 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_125
timestamp 1636968456
transform 1 0 12604 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_137
timestamp 1636968456
transform 1 0 13708 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_149
timestamp 1636968456
transform 1 0 14812 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_161
timestamp 1
transform 1 0 15916 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_167
timestamp 1
transform 1 0 16468 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_169
timestamp 1636968456
transform 1 0 16652 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_181
timestamp 1636968456
transform 1 0 17756 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_193
timestamp 1636968456
transform 1 0 18860 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_205
timestamp 1636968456
transform 1 0 19964 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_217
timestamp 1
transform 1 0 21068 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_223
timestamp 1
transform 1 0 21620 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_225
timestamp 1636968456
transform 1 0 21804 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_237
timestamp 1636968456
transform 1 0 22908 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_249
timestamp 1636968456
transform 1 0 24012 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_261
timestamp 1636968456
transform 1 0 25116 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_273
timestamp 1
transform 1 0 26220 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_279
timestamp 1
transform 1 0 26772 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_281
timestamp 1636968456
transform 1 0 26956 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_293
timestamp 1636968456
transform 1 0 28060 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_305
timestamp 1636968456
transform 1 0 29164 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_317
timestamp 1636968456
transform 1 0 30268 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_329
timestamp 1
transform 1 0 31372 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_335
timestamp 1
transform 1 0 31924 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_337
timestamp 1636968456
transform 1 0 32108 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_349
timestamp 1636968456
transform 1 0 33212 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_361
timestamp 1636968456
transform 1 0 34316 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_373
timestamp 1636968456
transform 1 0 35420 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_385
timestamp 1
transform 1 0 36524 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_391
timestamp 1
transform 1 0 37076 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_393
timestamp 1636968456
transform 1 0 37260 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_405
timestamp 1636968456
transform 1 0 38364 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_417
timestamp 1636968456
transform 1 0 39468 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_429
timestamp 1636968456
transform 1 0 40572 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_137_441
timestamp 1
transform 1 0 41676 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_137_444
timestamp 1
transform 1 0 41952 0 -1 77248
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_137_449
timestamp 1636968456
transform 1 0 42412 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_137_461
timestamp 1
transform 1 0 43516 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_137_482
timestamp 1
transform 1 0 45448 0 -1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_137_487
timestamp 1636968456
transform 1 0 45908 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_137_499
timestamp 1
transform 1 0 47012 0 -1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_137_503
timestamp 1
transform 1 0 47380 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_137_505
timestamp 1
transform 1 0 47564 0 -1 77248
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_137_511
timestamp 1636968456
transform 1 0 48116 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_137_523
timestamp 1
transform 1 0 49220 0 -1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_137_545
timestamp 1
transform 1 0 51244 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_548
timestamp 1636968456
transform 1 0 51520 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_561
timestamp 1
transform 1 0 52716 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_567
timestamp 1
transform 1 0 53268 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_570
timestamp 1636968456
transform 1 0 53544 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_137_582
timestamp 1
transform 1 0 54648 0 -1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_137_590
timestamp 1
transform 1 0 55384 0 -1 77248
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_137_594
timestamp 1636968456
transform 1 0 55752 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_606
timestamp 1
transform 1 0 56856 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_137_614
timestamp 1
transform 1 0 57592 0 -1 77248
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_137_617
timestamp 1636968456
transform 1 0 57868 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_629
timestamp 1636968456
transform 1 0 58972 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_641
timestamp 1636968456
transform 1 0 60076 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_653
timestamp 1636968456
transform 1 0 61180 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_665
timestamp 1
transform 1 0 62284 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_671
timestamp 1
transform 1 0 62836 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_673
timestamp 1636968456
transform 1 0 63020 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_685
timestamp 1636968456
transform 1 0 64124 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_697
timestamp 1636968456
transform 1 0 65228 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_709
timestamp 1636968456
transform 1 0 66332 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_721
timestamp 1
transform 1 0 67436 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_727
timestamp 1
transform 1 0 67988 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_729
timestamp 1636968456
transform 1 0 68172 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_741
timestamp 1636968456
transform 1 0 69276 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_753
timestamp 1636968456
transform 1 0 70380 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_765
timestamp 1636968456
transform 1 0 71484 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_777
timestamp 1
transform 1 0 72588 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_783
timestamp 1
transform 1 0 73140 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_785
timestamp 1636968456
transform 1 0 73324 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_797
timestamp 1636968456
transform 1 0 74428 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_809
timestamp 1636968456
transform 1 0 75532 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_821
timestamp 1636968456
transform 1 0 76636 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_833
timestamp 1
transform 1 0 77740 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_839
timestamp 1
transform 1 0 78292 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_841
timestamp 1636968456
transform 1 0 78476 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_853
timestamp 1636968456
transform 1 0 79580 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_865
timestamp 1636968456
transform 1 0 80684 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_877
timestamp 1636968456
transform 1 0 81788 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_889
timestamp 1
transform 1 0 82892 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_895
timestamp 1
transform 1 0 83444 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_897
timestamp 1636968456
transform 1 0 83628 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_909
timestamp 1636968456
transform 1 0 84732 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_921
timestamp 1636968456
transform 1 0 85836 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_933
timestamp 1636968456
transform 1 0 86940 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_945
timestamp 1
transform 1 0 88044 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_951
timestamp 1
transform 1 0 88596 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_953
timestamp 1636968456
transform 1 0 88780 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_965
timestamp 1636968456
transform 1 0 89884 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_977
timestamp 1636968456
transform 1 0 90988 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_989
timestamp 1636968456
transform 1 0 92092 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_1001
timestamp 1
transform 1 0 93196 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_1007
timestamp 1
transform 1 0 93748 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_1009
timestamp 1636968456
transform 1 0 93932 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_1021
timestamp 1636968456
transform 1 0 95036 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_1033
timestamp 1636968456
transform 1 0 96140 0 -1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_137_1045
timestamp 1636968456
transform 1 0 97244 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_137_1057
timestamp 1
transform 1 0 98348 0 -1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_1063
timestamp 1
transform 1 0 98900 0 -1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_1065
timestamp 1636968456
transform 1 0 99084 0 -1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_137_1077
timestamp 1
transform 1 0 100188 0 -1 77248
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_138_3
timestamp 1636968456
transform 1 0 1380 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_15
timestamp 1636968456
transform 1 0 2484 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_138_27
timestamp 1
transform 1 0 3588 0 1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_138_29
timestamp 1636968456
transform 1 0 3772 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_41
timestamp 1636968456
transform 1 0 4876 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_53
timestamp 1636968456
transform 1 0 5980 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_65
timestamp 1636968456
transform 1 0 7084 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_138_77
timestamp 1
transform 1 0 8188 0 1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_138_83
timestamp 1
transform 1 0 8740 0 1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_138_85
timestamp 1636968456
transform 1 0 8924 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_97
timestamp 1636968456
transform 1 0 10028 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_109
timestamp 1636968456
transform 1 0 11132 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_121
timestamp 1636968456
transform 1 0 12236 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_138_133
timestamp 1
transform 1 0 13340 0 1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_138_139
timestamp 1
transform 1 0 13892 0 1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_138_141
timestamp 1636968456
transform 1 0 14076 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_153
timestamp 1636968456
transform 1 0 15180 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_165
timestamp 1636968456
transform 1 0 16284 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_177
timestamp 1636968456
transform 1 0 17388 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_138_189
timestamp 1
transform 1 0 18492 0 1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_138_195
timestamp 1
transform 1 0 19044 0 1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_138_197
timestamp 1636968456
transform 1 0 19228 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_209
timestamp 1636968456
transform 1 0 20332 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_221
timestamp 1636968456
transform 1 0 21436 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_233
timestamp 1636968456
transform 1 0 22540 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_138_245
timestamp 1
transform 1 0 23644 0 1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_138_251
timestamp 1
transform 1 0 24196 0 1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_138_253
timestamp 1636968456
transform 1 0 24380 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_265
timestamp 1636968456
transform 1 0 25484 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_277
timestamp 1636968456
transform 1 0 26588 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_289
timestamp 1636968456
transform 1 0 27692 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_138_301
timestamp 1
transform 1 0 28796 0 1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_138_307
timestamp 1
transform 1 0 29348 0 1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_138_309
timestamp 1636968456
transform 1 0 29532 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_321
timestamp 1636968456
transform 1 0 30636 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_333
timestamp 1636968456
transform 1 0 31740 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_345
timestamp 1636968456
transform 1 0 32844 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_138_357
timestamp 1
transform 1 0 33948 0 1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_138_363
timestamp 1
transform 1 0 34500 0 1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_138_365
timestamp 1636968456
transform 1 0 34684 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_377
timestamp 1636968456
transform 1 0 35788 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_389
timestamp 1636968456
transform 1 0 36892 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_401
timestamp 1636968456
transform 1 0 37996 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_138_413
timestamp 1
transform 1 0 39100 0 1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_138_419
timestamp 1
transform 1 0 39652 0 1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_138_421
timestamp 1636968456
transform 1 0 39836 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_138_433
timestamp 1
transform 1 0 40940 0 1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_138_439
timestamp 1
transform 1 0 41492 0 1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_138_462
timestamp 1636968456
transform 1 0 43608 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_138_474
timestamp 1
transform 1 0 44712 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_138_477
timestamp 1
transform 1 0 44988 0 1 77248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_138_505
timestamp 1
transform 1 0 47564 0 1 77248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_138_529
timestamp 1
transform 1 0 49772 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_533
timestamp 1636968456
transform 1 0 50140 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_138_545
timestamp 1
transform 1 0 51244 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_138_566
timestamp 1
transform 1 0 53176 0 1 77248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_138_589
timestamp 1
transform 1 0 55292 0 1 77248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_138_632
timestamp 1636968456
transform 1 0 59248 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_645
timestamp 1636968456
transform 1 0 60444 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_657
timestamp 1636968456
transform 1 0 61548 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_669
timestamp 1636968456
transform 1 0 62652 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_681
timestamp 1636968456
transform 1 0 63756 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_138_693
timestamp 1
transform 1 0 64860 0 1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_138_699
timestamp 1
transform 1 0 65412 0 1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_138_701
timestamp 1636968456
transform 1 0 65596 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_713
timestamp 1636968456
transform 1 0 66700 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_725
timestamp 1636968456
transform 1 0 67804 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_737
timestamp 1636968456
transform 1 0 68908 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_138_749
timestamp 1
transform 1 0 70012 0 1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_138_755
timestamp 1
transform 1 0 70564 0 1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_138_757
timestamp 1636968456
transform 1 0 70748 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_769
timestamp 1636968456
transform 1 0 71852 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_781
timestamp 1636968456
transform 1 0 72956 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_793
timestamp 1636968456
transform 1 0 74060 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_138_805
timestamp 1
transform 1 0 75164 0 1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_138_811
timestamp 1
transform 1 0 75716 0 1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_138_813
timestamp 1636968456
transform 1 0 75900 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_825
timestamp 1636968456
transform 1 0 77004 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_837
timestamp 1636968456
transform 1 0 78108 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_849
timestamp 1636968456
transform 1 0 79212 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_138_861
timestamp 1
transform 1 0 80316 0 1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_138_867
timestamp 1
transform 1 0 80868 0 1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_138_869
timestamp 1636968456
transform 1 0 81052 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_881
timestamp 1636968456
transform 1 0 82156 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_893
timestamp 1636968456
transform 1 0 83260 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_905
timestamp 1636968456
transform 1 0 84364 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_138_917
timestamp 1
transform 1 0 85468 0 1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_138_923
timestamp 1
transform 1 0 86020 0 1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_138_925
timestamp 1636968456
transform 1 0 86204 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_937
timestamp 1636968456
transform 1 0 87308 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_949
timestamp 1636968456
transform 1 0 88412 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_961
timestamp 1636968456
transform 1 0 89516 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_138_973
timestamp 1
transform 1 0 90620 0 1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_138_979
timestamp 1
transform 1 0 91172 0 1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_138_981
timestamp 1636968456
transform 1 0 91356 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_993
timestamp 1636968456
transform 1 0 92460 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_1005
timestamp 1636968456
transform 1 0 93564 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_1017
timestamp 1636968456
transform 1 0 94668 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_138_1029
timestamp 1
transform 1 0 95772 0 1 77248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_138_1035
timestamp 1
transform 1 0 96324 0 1 77248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_138_1037
timestamp 1636968456
transform 1 0 96508 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_1049
timestamp 1636968456
transform 1 0 97612 0 1 77248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_1061
timestamp 1636968456
transform 1 0 98716 0 1 77248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_138_1073
timestamp 1
transform 1 0 99820 0 1 77248
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_139_3
timestamp 1636968456
transform 1 0 1380 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_15
timestamp 1636968456
transform 1 0 2484 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_27
timestamp 1636968456
transform 1 0 3588 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_39
timestamp 1636968456
transform 1 0 4692 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_139_51
timestamp 1
transform 1 0 5796 0 -1 78336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_139_55
timestamp 1
transform 1 0 6164 0 -1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_139_57
timestamp 1636968456
transform 1 0 6348 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_69
timestamp 1636968456
transform 1 0 7452 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_81
timestamp 1636968456
transform 1 0 8556 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_93
timestamp 1636968456
transform 1 0 9660 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_139_105
timestamp 1
transform 1 0 10764 0 -1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_139_111
timestamp 1
transform 1 0 11316 0 -1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_139_113
timestamp 1636968456
transform 1 0 11500 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_125
timestamp 1636968456
transform 1 0 12604 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_137
timestamp 1636968456
transform 1 0 13708 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_149
timestamp 1636968456
transform 1 0 14812 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_139_161
timestamp 1
transform 1 0 15916 0 -1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_139_167
timestamp 1
transform 1 0 16468 0 -1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_139_169
timestamp 1636968456
transform 1 0 16652 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_181
timestamp 1636968456
transform 1 0 17756 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_193
timestamp 1636968456
transform 1 0 18860 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_205
timestamp 1636968456
transform 1 0 19964 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_139_217
timestamp 1
transform 1 0 21068 0 -1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_139_223
timestamp 1
transform 1 0 21620 0 -1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_139_225
timestamp 1636968456
transform 1 0 21804 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_237
timestamp 1636968456
transform 1 0 22908 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_249
timestamp 1636968456
transform 1 0 24012 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_261
timestamp 1636968456
transform 1 0 25116 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_139_273
timestamp 1
transform 1 0 26220 0 -1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_139_279
timestamp 1
transform 1 0 26772 0 -1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_139_281
timestamp 1636968456
transform 1 0 26956 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_293
timestamp 1636968456
transform 1 0 28060 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_305
timestamp 1636968456
transform 1 0 29164 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_317
timestamp 1636968456
transform 1 0 30268 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_139_329
timestamp 1
transform 1 0 31372 0 -1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_139_335
timestamp 1
transform 1 0 31924 0 -1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_139_337
timestamp 1636968456
transform 1 0 32108 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_349
timestamp 1636968456
transform 1 0 33212 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_361
timestamp 1636968456
transform 1 0 34316 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_373
timestamp 1636968456
transform 1 0 35420 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_139_385
timestamp 1
transform 1 0 36524 0 -1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_139_391
timestamp 1
transform 1 0 37076 0 -1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_139_393
timestamp 1636968456
transform 1 0 37260 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_405
timestamp 1636968456
transform 1 0 38364 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_417
timestamp 1636968456
transform 1 0 39468 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_429
timestamp 1636968456
transform 1 0 40572 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_139_441
timestamp 1
transform 1 0 41676 0 -1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_139_447
timestamp 1
transform 1 0 42228 0 -1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_139_449
timestamp 1636968456
transform 1 0 42412 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_461
timestamp 1636968456
transform 1 0 43516 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_473
timestamp 1636968456
transform 1 0 44620 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_485
timestamp 1636968456
transform 1 0 45724 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_139_497
timestamp 1
transform 1 0 46828 0 -1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_139_503
timestamp 1
transform 1 0 47380 0 -1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_139_505
timestamp 1636968456
transform 1 0 47564 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_517
timestamp 1636968456
transform 1 0 48668 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_529
timestamp 1636968456
transform 1 0 49772 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_541
timestamp 1636968456
transform 1 0 50876 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_139_553
timestamp 1
transform 1 0 51980 0 -1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_139_559
timestamp 1
transform 1 0 52532 0 -1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_139_561
timestamp 1636968456
transform 1 0 52716 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_573
timestamp 1636968456
transform 1 0 53820 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_585
timestamp 1636968456
transform 1 0 54924 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_597
timestamp 1636968456
transform 1 0 56028 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_139_609
timestamp 1
transform 1 0 57132 0 -1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_139_615
timestamp 1
transform 1 0 57684 0 -1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_139_617
timestamp 1636968456
transform 1 0 57868 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_629
timestamp 1636968456
transform 1 0 58972 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_641
timestamp 1636968456
transform 1 0 60076 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_653
timestamp 1636968456
transform 1 0 61180 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_139_665
timestamp 1
transform 1 0 62284 0 -1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_139_671
timestamp 1
transform 1 0 62836 0 -1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_139_673
timestamp 1636968456
transform 1 0 63020 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_685
timestamp 1636968456
transform 1 0 64124 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_697
timestamp 1636968456
transform 1 0 65228 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_709
timestamp 1636968456
transform 1 0 66332 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_139_721
timestamp 1
transform 1 0 67436 0 -1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_139_727
timestamp 1
transform 1 0 67988 0 -1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_139_729
timestamp 1636968456
transform 1 0 68172 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_741
timestamp 1636968456
transform 1 0 69276 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_753
timestamp 1636968456
transform 1 0 70380 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_765
timestamp 1636968456
transform 1 0 71484 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_139_777
timestamp 1
transform 1 0 72588 0 -1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_139_783
timestamp 1
transform 1 0 73140 0 -1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_139_785
timestamp 1636968456
transform 1 0 73324 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_797
timestamp 1636968456
transform 1 0 74428 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_809
timestamp 1636968456
transform 1 0 75532 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_821
timestamp 1636968456
transform 1 0 76636 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_139_833
timestamp 1
transform 1 0 77740 0 -1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_139_839
timestamp 1
transform 1 0 78292 0 -1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_139_841
timestamp 1636968456
transform 1 0 78476 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_853
timestamp 1636968456
transform 1 0 79580 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_865
timestamp 1636968456
transform 1 0 80684 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_877
timestamp 1636968456
transform 1 0 81788 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_139_889
timestamp 1
transform 1 0 82892 0 -1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_139_895
timestamp 1
transform 1 0 83444 0 -1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_139_897
timestamp 1636968456
transform 1 0 83628 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_909
timestamp 1636968456
transform 1 0 84732 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_921
timestamp 1636968456
transform 1 0 85836 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_933
timestamp 1636968456
transform 1 0 86940 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_139_945
timestamp 1
transform 1 0 88044 0 -1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_139_951
timestamp 1
transform 1 0 88596 0 -1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_139_953
timestamp 1636968456
transform 1 0 88780 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_965
timestamp 1636968456
transform 1 0 89884 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_977
timestamp 1636968456
transform 1 0 90988 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_989
timestamp 1636968456
transform 1 0 92092 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_139_1001
timestamp 1
transform 1 0 93196 0 -1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_139_1007
timestamp 1
transform 1 0 93748 0 -1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_139_1009
timestamp 1636968456
transform 1 0 93932 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_1021
timestamp 1636968456
transform 1 0 95036 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_1033
timestamp 1636968456
transform 1 0 96140 0 -1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_139_1045
timestamp 1636968456
transform 1 0 97244 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_139_1057
timestamp 1
transform 1 0 98348 0 -1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_139_1063
timestamp 1
transform 1 0 98900 0 -1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_139_1065
timestamp 1636968456
transform 1 0 99084 0 -1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_139_1077
timestamp 1
transform 1 0 100188 0 -1 78336
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_140_3
timestamp 1636968456
transform 1 0 1380 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_15
timestamp 1636968456
transform 1 0 2484 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_140_27
timestamp 1
transform 1 0 3588 0 1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_140_29
timestamp 1636968456
transform 1 0 3772 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_41
timestamp 1636968456
transform 1 0 4876 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_53
timestamp 1636968456
transform 1 0 5980 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_65
timestamp 1636968456
transform 1 0 7084 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_140_77
timestamp 1
transform 1 0 8188 0 1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_140_83
timestamp 1
transform 1 0 8740 0 1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_140_85
timestamp 1636968456
transform 1 0 8924 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_97
timestamp 1636968456
transform 1 0 10028 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_109
timestamp 1636968456
transform 1 0 11132 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_121
timestamp 1636968456
transform 1 0 12236 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_140_133
timestamp 1
transform 1 0 13340 0 1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_140_139
timestamp 1
transform 1 0 13892 0 1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_140_141
timestamp 1636968456
transform 1 0 14076 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_153
timestamp 1636968456
transform 1 0 15180 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_165
timestamp 1636968456
transform 1 0 16284 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_177
timestamp 1636968456
transform 1 0 17388 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_140_189
timestamp 1
transform 1 0 18492 0 1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_140_195
timestamp 1
transform 1 0 19044 0 1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_140_197
timestamp 1636968456
transform 1 0 19228 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_209
timestamp 1636968456
transform 1 0 20332 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_221
timestamp 1636968456
transform 1 0 21436 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_233
timestamp 1636968456
transform 1 0 22540 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_140_245
timestamp 1
transform 1 0 23644 0 1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_140_251
timestamp 1
transform 1 0 24196 0 1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_140_253
timestamp 1636968456
transform 1 0 24380 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_265
timestamp 1636968456
transform 1 0 25484 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_277
timestamp 1636968456
transform 1 0 26588 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_289
timestamp 1636968456
transform 1 0 27692 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_140_301
timestamp 1
transform 1 0 28796 0 1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_140_307
timestamp 1
transform 1 0 29348 0 1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_140_309
timestamp 1636968456
transform 1 0 29532 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_321
timestamp 1636968456
transform 1 0 30636 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_333
timestamp 1636968456
transform 1 0 31740 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_345
timestamp 1636968456
transform 1 0 32844 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_140_357
timestamp 1
transform 1 0 33948 0 1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_140_363
timestamp 1
transform 1 0 34500 0 1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_140_365
timestamp 1636968456
transform 1 0 34684 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_377
timestamp 1636968456
transform 1 0 35788 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_389
timestamp 1636968456
transform 1 0 36892 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_401
timestamp 1636968456
transform 1 0 37996 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_140_413
timestamp 1
transform 1 0 39100 0 1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_140_419
timestamp 1
transform 1 0 39652 0 1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_140_421
timestamp 1636968456
transform 1 0 39836 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_433
timestamp 1636968456
transform 1 0 40940 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_445
timestamp 1636968456
transform 1 0 42044 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_457
timestamp 1636968456
transform 1 0 43148 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_140_469
timestamp 1
transform 1 0 44252 0 1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_140_475
timestamp 1
transform 1 0 44804 0 1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_140_477
timestamp 1636968456
transform 1 0 44988 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_489
timestamp 1636968456
transform 1 0 46092 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_501
timestamp 1636968456
transform 1 0 47196 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_513
timestamp 1636968456
transform 1 0 48300 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_140_525
timestamp 1
transform 1 0 49404 0 1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_140_531
timestamp 1
transform 1 0 49956 0 1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_140_533
timestamp 1636968456
transform 1 0 50140 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_545
timestamp 1636968456
transform 1 0 51244 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_557
timestamp 1636968456
transform 1 0 52348 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_569
timestamp 1636968456
transform 1 0 53452 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_140_581
timestamp 1
transform 1 0 54556 0 1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_140_587
timestamp 1
transform 1 0 55108 0 1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_140_589
timestamp 1636968456
transform 1 0 55292 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_601
timestamp 1636968456
transform 1 0 56396 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_613
timestamp 1636968456
transform 1 0 57500 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_625
timestamp 1636968456
transform 1 0 58604 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_140_637
timestamp 1
transform 1 0 59708 0 1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_140_643
timestamp 1
transform 1 0 60260 0 1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_140_645
timestamp 1636968456
transform 1 0 60444 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_657
timestamp 1636968456
transform 1 0 61548 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_669
timestamp 1636968456
transform 1 0 62652 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_681
timestamp 1636968456
transform 1 0 63756 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_140_693
timestamp 1
transform 1 0 64860 0 1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_140_699
timestamp 1
transform 1 0 65412 0 1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_140_701
timestamp 1636968456
transform 1 0 65596 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_713
timestamp 1636968456
transform 1 0 66700 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_725
timestamp 1636968456
transform 1 0 67804 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_737
timestamp 1636968456
transform 1 0 68908 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_140_749
timestamp 1
transform 1 0 70012 0 1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_140_755
timestamp 1
transform 1 0 70564 0 1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_140_757
timestamp 1636968456
transform 1 0 70748 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_769
timestamp 1636968456
transform 1 0 71852 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_781
timestamp 1636968456
transform 1 0 72956 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_793
timestamp 1636968456
transform 1 0 74060 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_140_805
timestamp 1
transform 1 0 75164 0 1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_140_811
timestamp 1
transform 1 0 75716 0 1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_140_813
timestamp 1636968456
transform 1 0 75900 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_825
timestamp 1636968456
transform 1 0 77004 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_837
timestamp 1636968456
transform 1 0 78108 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_849
timestamp 1636968456
transform 1 0 79212 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_140_861
timestamp 1
transform 1 0 80316 0 1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_140_867
timestamp 1
transform 1 0 80868 0 1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_140_869
timestamp 1636968456
transform 1 0 81052 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_881
timestamp 1636968456
transform 1 0 82156 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_893
timestamp 1636968456
transform 1 0 83260 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_905
timestamp 1636968456
transform 1 0 84364 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_140_917
timestamp 1
transform 1 0 85468 0 1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_140_923
timestamp 1
transform 1 0 86020 0 1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_140_925
timestamp 1636968456
transform 1 0 86204 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_937
timestamp 1636968456
transform 1 0 87308 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_949
timestamp 1636968456
transform 1 0 88412 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_961
timestamp 1636968456
transform 1 0 89516 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_140_973
timestamp 1
transform 1 0 90620 0 1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_140_979
timestamp 1
transform 1 0 91172 0 1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_140_981
timestamp 1636968456
transform 1 0 91356 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_993
timestamp 1636968456
transform 1 0 92460 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_1005
timestamp 1636968456
transform 1 0 93564 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_1017
timestamp 1636968456
transform 1 0 94668 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_140_1029
timestamp 1
transform 1 0 95772 0 1 78336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_140_1035
timestamp 1
transform 1 0 96324 0 1 78336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_140_1037
timestamp 1636968456
transform 1 0 96508 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_1049
timestamp 1636968456
transform 1 0 97612 0 1 78336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_1061
timestamp 1636968456
transform 1 0 98716 0 1 78336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_140_1073
timestamp 1
transform 1 0 99820 0 1 78336
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_141_3
timestamp 1636968456
transform 1 0 1380 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_15
timestamp 1636968456
transform 1 0 2484 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_27
timestamp 1636968456
transform 1 0 3588 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_39
timestamp 1636968456
transform 1 0 4692 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_141_51
timestamp 1
transform 1 0 5796 0 -1 79424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_141_55
timestamp 1
transform 1 0 6164 0 -1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_141_57
timestamp 1636968456
transform 1 0 6348 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_69
timestamp 1636968456
transform 1 0 7452 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_81
timestamp 1636968456
transform 1 0 8556 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_93
timestamp 1636968456
transform 1 0 9660 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_141_105
timestamp 1
transform 1 0 10764 0 -1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_141_111
timestamp 1
transform 1 0 11316 0 -1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_141_113
timestamp 1636968456
transform 1 0 11500 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_125
timestamp 1636968456
transform 1 0 12604 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_137
timestamp 1636968456
transform 1 0 13708 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_149
timestamp 1636968456
transform 1 0 14812 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_141_161
timestamp 1
transform 1 0 15916 0 -1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_141_167
timestamp 1
transform 1 0 16468 0 -1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_141_169
timestamp 1636968456
transform 1 0 16652 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_181
timestamp 1636968456
transform 1 0 17756 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_193
timestamp 1636968456
transform 1 0 18860 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_205
timestamp 1636968456
transform 1 0 19964 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_141_217
timestamp 1
transform 1 0 21068 0 -1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_141_223
timestamp 1
transform 1 0 21620 0 -1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_141_225
timestamp 1636968456
transform 1 0 21804 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_237
timestamp 1636968456
transform 1 0 22908 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_249
timestamp 1636968456
transform 1 0 24012 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_261
timestamp 1636968456
transform 1 0 25116 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_141_273
timestamp 1
transform 1 0 26220 0 -1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_141_279
timestamp 1
transform 1 0 26772 0 -1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_141_281
timestamp 1636968456
transform 1 0 26956 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_293
timestamp 1636968456
transform 1 0 28060 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_305
timestamp 1636968456
transform 1 0 29164 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_317
timestamp 1636968456
transform 1 0 30268 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_141_329
timestamp 1
transform 1 0 31372 0 -1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_141_335
timestamp 1
transform 1 0 31924 0 -1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_141_337
timestamp 1636968456
transform 1 0 32108 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_349
timestamp 1636968456
transform 1 0 33212 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_361
timestamp 1636968456
transform 1 0 34316 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_373
timestamp 1636968456
transform 1 0 35420 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_141_385
timestamp 1
transform 1 0 36524 0 -1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_141_391
timestamp 1
transform 1 0 37076 0 -1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_141_393
timestamp 1636968456
transform 1 0 37260 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_405
timestamp 1636968456
transform 1 0 38364 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_417
timestamp 1636968456
transform 1 0 39468 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_429
timestamp 1636968456
transform 1 0 40572 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_141_441
timestamp 1
transform 1 0 41676 0 -1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_141_447
timestamp 1
transform 1 0 42228 0 -1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_141_449
timestamp 1636968456
transform 1 0 42412 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_461
timestamp 1636968456
transform 1 0 43516 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_473
timestamp 1636968456
transform 1 0 44620 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_485
timestamp 1636968456
transform 1 0 45724 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_141_497
timestamp 1
transform 1 0 46828 0 -1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_141_503
timestamp 1
transform 1 0 47380 0 -1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_141_505
timestamp 1636968456
transform 1 0 47564 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_517
timestamp 1636968456
transform 1 0 48668 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_529
timestamp 1636968456
transform 1 0 49772 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_541
timestamp 1636968456
transform 1 0 50876 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_141_553
timestamp 1
transform 1 0 51980 0 -1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_141_559
timestamp 1
transform 1 0 52532 0 -1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_141_561
timestamp 1636968456
transform 1 0 52716 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_573
timestamp 1636968456
transform 1 0 53820 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_585
timestamp 1636968456
transform 1 0 54924 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_597
timestamp 1636968456
transform 1 0 56028 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_141_609
timestamp 1
transform 1 0 57132 0 -1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_141_615
timestamp 1
transform 1 0 57684 0 -1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_141_617
timestamp 1636968456
transform 1 0 57868 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_629
timestamp 1636968456
transform 1 0 58972 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_641
timestamp 1636968456
transform 1 0 60076 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_653
timestamp 1636968456
transform 1 0 61180 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_141_665
timestamp 1
transform 1 0 62284 0 -1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_141_671
timestamp 1
transform 1 0 62836 0 -1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_141_673
timestamp 1636968456
transform 1 0 63020 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_685
timestamp 1636968456
transform 1 0 64124 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_697
timestamp 1636968456
transform 1 0 65228 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_709
timestamp 1636968456
transform 1 0 66332 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_141_721
timestamp 1
transform 1 0 67436 0 -1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_141_727
timestamp 1
transform 1 0 67988 0 -1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_141_729
timestamp 1636968456
transform 1 0 68172 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_741
timestamp 1636968456
transform 1 0 69276 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_753
timestamp 1636968456
transform 1 0 70380 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_765
timestamp 1636968456
transform 1 0 71484 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_141_777
timestamp 1
transform 1 0 72588 0 -1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_141_783
timestamp 1
transform 1 0 73140 0 -1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_141_785
timestamp 1636968456
transform 1 0 73324 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_797
timestamp 1636968456
transform 1 0 74428 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_809
timestamp 1636968456
transform 1 0 75532 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_821
timestamp 1636968456
transform 1 0 76636 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_141_833
timestamp 1
transform 1 0 77740 0 -1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_141_839
timestamp 1
transform 1 0 78292 0 -1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_141_841
timestamp 1636968456
transform 1 0 78476 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_853
timestamp 1636968456
transform 1 0 79580 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_865
timestamp 1636968456
transform 1 0 80684 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_877
timestamp 1636968456
transform 1 0 81788 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_141_889
timestamp 1
transform 1 0 82892 0 -1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_141_895
timestamp 1
transform 1 0 83444 0 -1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_141_897
timestamp 1636968456
transform 1 0 83628 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_909
timestamp 1636968456
transform 1 0 84732 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_921
timestamp 1636968456
transform 1 0 85836 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_933
timestamp 1636968456
transform 1 0 86940 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_141_945
timestamp 1
transform 1 0 88044 0 -1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_141_951
timestamp 1
transform 1 0 88596 0 -1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_141_953
timestamp 1636968456
transform 1 0 88780 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_965
timestamp 1636968456
transform 1 0 89884 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_977
timestamp 1636968456
transform 1 0 90988 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_989
timestamp 1636968456
transform 1 0 92092 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_141_1001
timestamp 1
transform 1 0 93196 0 -1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_141_1007
timestamp 1
transform 1 0 93748 0 -1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_141_1009
timestamp 1636968456
transform 1 0 93932 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_1021
timestamp 1636968456
transform 1 0 95036 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_1033
timestamp 1636968456
transform 1 0 96140 0 -1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_1045
timestamp 1636968456
transform 1 0 97244 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_141_1057
timestamp 1
transform 1 0 98348 0 -1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_141_1063
timestamp 1
transform 1 0 98900 0 -1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_141_1065
timestamp 1636968456
transform 1 0 99084 0 -1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_141_1077
timestamp 1
transform 1 0 100188 0 -1 79424
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_142_3
timestamp 1636968456
transform 1 0 1380 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_15
timestamp 1636968456
transform 1 0 2484 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_142_27
timestamp 1
transform 1 0 3588 0 1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_142_29
timestamp 1636968456
transform 1 0 3772 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_41
timestamp 1636968456
transform 1 0 4876 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_53
timestamp 1636968456
transform 1 0 5980 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_65
timestamp 1636968456
transform 1 0 7084 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_142_77
timestamp 1
transform 1 0 8188 0 1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_142_83
timestamp 1
transform 1 0 8740 0 1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_142_85
timestamp 1636968456
transform 1 0 8924 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_97
timestamp 1636968456
transform 1 0 10028 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_109
timestamp 1636968456
transform 1 0 11132 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_121
timestamp 1636968456
transform 1 0 12236 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_142_133
timestamp 1
transform 1 0 13340 0 1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_142_139
timestamp 1
transform 1 0 13892 0 1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_142_141
timestamp 1636968456
transform 1 0 14076 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_153
timestamp 1636968456
transform 1 0 15180 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_165
timestamp 1636968456
transform 1 0 16284 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_177
timestamp 1636968456
transform 1 0 17388 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_142_189
timestamp 1
transform 1 0 18492 0 1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_142_195
timestamp 1
transform 1 0 19044 0 1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_142_197
timestamp 1636968456
transform 1 0 19228 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_209
timestamp 1636968456
transform 1 0 20332 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_221
timestamp 1636968456
transform 1 0 21436 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_233
timestamp 1636968456
transform 1 0 22540 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_142_245
timestamp 1
transform 1 0 23644 0 1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_142_251
timestamp 1
transform 1 0 24196 0 1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_142_253
timestamp 1636968456
transform 1 0 24380 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_265
timestamp 1636968456
transform 1 0 25484 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_277
timestamp 1636968456
transform 1 0 26588 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_289
timestamp 1636968456
transform 1 0 27692 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_142_301
timestamp 1
transform 1 0 28796 0 1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_142_307
timestamp 1
transform 1 0 29348 0 1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_142_309
timestamp 1636968456
transform 1 0 29532 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_321
timestamp 1636968456
transform 1 0 30636 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_333
timestamp 1636968456
transform 1 0 31740 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_345
timestamp 1636968456
transform 1 0 32844 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_142_357
timestamp 1
transform 1 0 33948 0 1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_142_363
timestamp 1
transform 1 0 34500 0 1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_142_365
timestamp 1636968456
transform 1 0 34684 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_377
timestamp 1636968456
transform 1 0 35788 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_389
timestamp 1636968456
transform 1 0 36892 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_401
timestamp 1636968456
transform 1 0 37996 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_142_413
timestamp 1
transform 1 0 39100 0 1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_142_419
timestamp 1
transform 1 0 39652 0 1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_142_421
timestamp 1636968456
transform 1 0 39836 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_433
timestamp 1636968456
transform 1 0 40940 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_445
timestamp 1636968456
transform 1 0 42044 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_457
timestamp 1636968456
transform 1 0 43148 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_142_469
timestamp 1
transform 1 0 44252 0 1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_142_475
timestamp 1
transform 1 0 44804 0 1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_142_477
timestamp 1636968456
transform 1 0 44988 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_489
timestamp 1636968456
transform 1 0 46092 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_501
timestamp 1636968456
transform 1 0 47196 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_513
timestamp 1636968456
transform 1 0 48300 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_142_525
timestamp 1
transform 1 0 49404 0 1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_142_531
timestamp 1
transform 1 0 49956 0 1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_142_533
timestamp 1636968456
transform 1 0 50140 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_545
timestamp 1636968456
transform 1 0 51244 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_557
timestamp 1636968456
transform 1 0 52348 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_569
timestamp 1636968456
transform 1 0 53452 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_142_581
timestamp 1
transform 1 0 54556 0 1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_142_587
timestamp 1
transform 1 0 55108 0 1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_142_589
timestamp 1636968456
transform 1 0 55292 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_601
timestamp 1636968456
transform 1 0 56396 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_613
timestamp 1636968456
transform 1 0 57500 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_625
timestamp 1636968456
transform 1 0 58604 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_142_637
timestamp 1
transform 1 0 59708 0 1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_142_643
timestamp 1
transform 1 0 60260 0 1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_142_645
timestamp 1636968456
transform 1 0 60444 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_657
timestamp 1636968456
transform 1 0 61548 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_669
timestamp 1636968456
transform 1 0 62652 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_681
timestamp 1636968456
transform 1 0 63756 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_142_693
timestamp 1
transform 1 0 64860 0 1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_142_699
timestamp 1
transform 1 0 65412 0 1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_142_701
timestamp 1636968456
transform 1 0 65596 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_713
timestamp 1636968456
transform 1 0 66700 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_725
timestamp 1636968456
transform 1 0 67804 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_737
timestamp 1636968456
transform 1 0 68908 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_142_749
timestamp 1
transform 1 0 70012 0 1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_142_755
timestamp 1
transform 1 0 70564 0 1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_142_757
timestamp 1636968456
transform 1 0 70748 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_769
timestamp 1636968456
transform 1 0 71852 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_781
timestamp 1636968456
transform 1 0 72956 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_793
timestamp 1636968456
transform 1 0 74060 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_142_805
timestamp 1
transform 1 0 75164 0 1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_142_811
timestamp 1
transform 1 0 75716 0 1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_142_813
timestamp 1636968456
transform 1 0 75900 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_825
timestamp 1636968456
transform 1 0 77004 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_837
timestamp 1636968456
transform 1 0 78108 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_849
timestamp 1636968456
transform 1 0 79212 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_142_861
timestamp 1
transform 1 0 80316 0 1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_142_867
timestamp 1
transform 1 0 80868 0 1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_142_869
timestamp 1636968456
transform 1 0 81052 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_881
timestamp 1636968456
transform 1 0 82156 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_893
timestamp 1636968456
transform 1 0 83260 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_905
timestamp 1636968456
transform 1 0 84364 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_142_917
timestamp 1
transform 1 0 85468 0 1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_142_923
timestamp 1
transform 1 0 86020 0 1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_142_925
timestamp 1636968456
transform 1 0 86204 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_937
timestamp 1636968456
transform 1 0 87308 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_949
timestamp 1636968456
transform 1 0 88412 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_961
timestamp 1636968456
transform 1 0 89516 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_142_973
timestamp 1
transform 1 0 90620 0 1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_142_979
timestamp 1
transform 1 0 91172 0 1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_142_981
timestamp 1636968456
transform 1 0 91356 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_993
timestamp 1636968456
transform 1 0 92460 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_1005
timestamp 1636968456
transform 1 0 93564 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_1017
timestamp 1636968456
transform 1 0 94668 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_142_1029
timestamp 1
transform 1 0 95772 0 1 79424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_142_1035
timestamp 1
transform 1 0 96324 0 1 79424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_142_1037
timestamp 1636968456
transform 1 0 96508 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_1049
timestamp 1636968456
transform 1 0 97612 0 1 79424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_1061
timestamp 1636968456
transform 1 0 98716 0 1 79424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_142_1073
timestamp 1
transform 1 0 99820 0 1 79424
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_143_3
timestamp 1636968456
transform 1 0 1380 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_15
timestamp 1636968456
transform 1 0 2484 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_27
timestamp 1636968456
transform 1 0 3588 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_39
timestamp 1636968456
transform 1 0 4692 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_143_51
timestamp 1
transform 1 0 5796 0 -1 80512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_143_55
timestamp 1
transform 1 0 6164 0 -1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_143_57
timestamp 1636968456
transform 1 0 6348 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_69
timestamp 1636968456
transform 1 0 7452 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_81
timestamp 1636968456
transform 1 0 8556 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_93
timestamp 1636968456
transform 1 0 9660 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_143_105
timestamp 1
transform 1 0 10764 0 -1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_143_111
timestamp 1
transform 1 0 11316 0 -1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_143_113
timestamp 1636968456
transform 1 0 11500 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_125
timestamp 1636968456
transform 1 0 12604 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_137
timestamp 1636968456
transform 1 0 13708 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_149
timestamp 1636968456
transform 1 0 14812 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_143_161
timestamp 1
transform 1 0 15916 0 -1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_143_167
timestamp 1
transform 1 0 16468 0 -1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_143_169
timestamp 1636968456
transform 1 0 16652 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_181
timestamp 1636968456
transform 1 0 17756 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_193
timestamp 1636968456
transform 1 0 18860 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_205
timestamp 1636968456
transform 1 0 19964 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_143_217
timestamp 1
transform 1 0 21068 0 -1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_143_223
timestamp 1
transform 1 0 21620 0 -1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_143_225
timestamp 1636968456
transform 1 0 21804 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_237
timestamp 1636968456
transform 1 0 22908 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_249
timestamp 1636968456
transform 1 0 24012 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_261
timestamp 1636968456
transform 1 0 25116 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_143_273
timestamp 1
transform 1 0 26220 0 -1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_143_279
timestamp 1
transform 1 0 26772 0 -1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_143_281
timestamp 1636968456
transform 1 0 26956 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_293
timestamp 1636968456
transform 1 0 28060 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_305
timestamp 1636968456
transform 1 0 29164 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_317
timestamp 1636968456
transform 1 0 30268 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_143_329
timestamp 1
transform 1 0 31372 0 -1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_143_335
timestamp 1
transform 1 0 31924 0 -1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_143_337
timestamp 1636968456
transform 1 0 32108 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_349
timestamp 1636968456
transform 1 0 33212 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_361
timestamp 1636968456
transform 1 0 34316 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_373
timestamp 1636968456
transform 1 0 35420 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_143_385
timestamp 1
transform 1 0 36524 0 -1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_143_391
timestamp 1
transform 1 0 37076 0 -1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_143_393
timestamp 1636968456
transform 1 0 37260 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_405
timestamp 1636968456
transform 1 0 38364 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_417
timestamp 1636968456
transform 1 0 39468 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_429
timestamp 1636968456
transform 1 0 40572 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_143_441
timestamp 1
transform 1 0 41676 0 -1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_143_447
timestamp 1
transform 1 0 42228 0 -1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_143_449
timestamp 1636968456
transform 1 0 42412 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_461
timestamp 1636968456
transform 1 0 43516 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_473
timestamp 1636968456
transform 1 0 44620 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_485
timestamp 1636968456
transform 1 0 45724 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_143_497
timestamp 1
transform 1 0 46828 0 -1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_143_503
timestamp 1
transform 1 0 47380 0 -1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_143_505
timestamp 1636968456
transform 1 0 47564 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_517
timestamp 1636968456
transform 1 0 48668 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_529
timestamp 1636968456
transform 1 0 49772 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_541
timestamp 1636968456
transform 1 0 50876 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_143_553
timestamp 1
transform 1 0 51980 0 -1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_143_559
timestamp 1
transform 1 0 52532 0 -1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_143_561
timestamp 1636968456
transform 1 0 52716 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_573
timestamp 1636968456
transform 1 0 53820 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_585
timestamp 1636968456
transform 1 0 54924 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_597
timestamp 1636968456
transform 1 0 56028 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_143_609
timestamp 1
transform 1 0 57132 0 -1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_143_615
timestamp 1
transform 1 0 57684 0 -1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_143_617
timestamp 1636968456
transform 1 0 57868 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_629
timestamp 1636968456
transform 1 0 58972 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_641
timestamp 1636968456
transform 1 0 60076 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_653
timestamp 1636968456
transform 1 0 61180 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_143_665
timestamp 1
transform 1 0 62284 0 -1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_143_671
timestamp 1
transform 1 0 62836 0 -1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_143_673
timestamp 1636968456
transform 1 0 63020 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_685
timestamp 1636968456
transform 1 0 64124 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_697
timestamp 1636968456
transform 1 0 65228 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_709
timestamp 1636968456
transform 1 0 66332 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_143_721
timestamp 1
transform 1 0 67436 0 -1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_143_727
timestamp 1
transform 1 0 67988 0 -1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_143_729
timestamp 1636968456
transform 1 0 68172 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_741
timestamp 1636968456
transform 1 0 69276 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_753
timestamp 1636968456
transform 1 0 70380 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_765
timestamp 1636968456
transform 1 0 71484 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_143_777
timestamp 1
transform 1 0 72588 0 -1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_143_783
timestamp 1
transform 1 0 73140 0 -1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_143_785
timestamp 1636968456
transform 1 0 73324 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_797
timestamp 1636968456
transform 1 0 74428 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_809
timestamp 1636968456
transform 1 0 75532 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_821
timestamp 1636968456
transform 1 0 76636 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_143_833
timestamp 1
transform 1 0 77740 0 -1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_143_839
timestamp 1
transform 1 0 78292 0 -1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_143_841
timestamp 1636968456
transform 1 0 78476 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_853
timestamp 1636968456
transform 1 0 79580 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_865
timestamp 1636968456
transform 1 0 80684 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_877
timestamp 1636968456
transform 1 0 81788 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_143_889
timestamp 1
transform 1 0 82892 0 -1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_143_895
timestamp 1
transform 1 0 83444 0 -1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_143_897
timestamp 1636968456
transform 1 0 83628 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_909
timestamp 1636968456
transform 1 0 84732 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_921
timestamp 1636968456
transform 1 0 85836 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_933
timestamp 1636968456
transform 1 0 86940 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_143_945
timestamp 1
transform 1 0 88044 0 -1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_143_951
timestamp 1
transform 1 0 88596 0 -1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_143_953
timestamp 1636968456
transform 1 0 88780 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_965
timestamp 1636968456
transform 1 0 89884 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_977
timestamp 1636968456
transform 1 0 90988 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_989
timestamp 1636968456
transform 1 0 92092 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_143_1001
timestamp 1
transform 1 0 93196 0 -1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_143_1007
timestamp 1
transform 1 0 93748 0 -1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_143_1009
timestamp 1636968456
transform 1 0 93932 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_1021
timestamp 1636968456
transform 1 0 95036 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_1033
timestamp 1636968456
transform 1 0 96140 0 -1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_1045
timestamp 1636968456
transform 1 0 97244 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_143_1057
timestamp 1
transform 1 0 98348 0 -1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_143_1063
timestamp 1
transform 1 0 98900 0 -1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_143_1065
timestamp 1636968456
transform 1 0 99084 0 -1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_143_1077
timestamp 1
transform 1 0 100188 0 -1 80512
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_144_3
timestamp 1636968456
transform 1 0 1380 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_15
timestamp 1636968456
transform 1 0 2484 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_144_27
timestamp 1
transform 1 0 3588 0 1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_144_29
timestamp 1636968456
transform 1 0 3772 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_41
timestamp 1636968456
transform 1 0 4876 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_53
timestamp 1636968456
transform 1 0 5980 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_65
timestamp 1636968456
transform 1 0 7084 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_144_77
timestamp 1
transform 1 0 8188 0 1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_144_83
timestamp 1
transform 1 0 8740 0 1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_144_85
timestamp 1636968456
transform 1 0 8924 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_97
timestamp 1636968456
transform 1 0 10028 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_109
timestamp 1636968456
transform 1 0 11132 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_121
timestamp 1636968456
transform 1 0 12236 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_144_133
timestamp 1
transform 1 0 13340 0 1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_144_139
timestamp 1
transform 1 0 13892 0 1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_144_141
timestamp 1636968456
transform 1 0 14076 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_153
timestamp 1636968456
transform 1 0 15180 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_165
timestamp 1636968456
transform 1 0 16284 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_177
timestamp 1636968456
transform 1 0 17388 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_144_189
timestamp 1
transform 1 0 18492 0 1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_144_195
timestamp 1
transform 1 0 19044 0 1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_144_197
timestamp 1636968456
transform 1 0 19228 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_209
timestamp 1636968456
transform 1 0 20332 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_221
timestamp 1636968456
transform 1 0 21436 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_233
timestamp 1636968456
transform 1 0 22540 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_144_245
timestamp 1
transform 1 0 23644 0 1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_144_251
timestamp 1
transform 1 0 24196 0 1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_144_253
timestamp 1636968456
transform 1 0 24380 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_265
timestamp 1636968456
transform 1 0 25484 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_277
timestamp 1636968456
transform 1 0 26588 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_289
timestamp 1636968456
transform 1 0 27692 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_144_301
timestamp 1
transform 1 0 28796 0 1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_144_307
timestamp 1
transform 1 0 29348 0 1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_144_309
timestamp 1636968456
transform 1 0 29532 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_321
timestamp 1636968456
transform 1 0 30636 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_333
timestamp 1636968456
transform 1 0 31740 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_345
timestamp 1636968456
transform 1 0 32844 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_144_357
timestamp 1
transform 1 0 33948 0 1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_144_363
timestamp 1
transform 1 0 34500 0 1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_144_365
timestamp 1636968456
transform 1 0 34684 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_377
timestamp 1636968456
transform 1 0 35788 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_389
timestamp 1636968456
transform 1 0 36892 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_401
timestamp 1636968456
transform 1 0 37996 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_144_413
timestamp 1
transform 1 0 39100 0 1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_144_419
timestamp 1
transform 1 0 39652 0 1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_144_421
timestamp 1636968456
transform 1 0 39836 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_433
timestamp 1636968456
transform 1 0 40940 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_445
timestamp 1636968456
transform 1 0 42044 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_457
timestamp 1636968456
transform 1 0 43148 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_144_469
timestamp 1
transform 1 0 44252 0 1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_144_475
timestamp 1
transform 1 0 44804 0 1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_144_477
timestamp 1636968456
transform 1 0 44988 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_489
timestamp 1636968456
transform 1 0 46092 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_501
timestamp 1636968456
transform 1 0 47196 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_513
timestamp 1636968456
transform 1 0 48300 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_144_525
timestamp 1
transform 1 0 49404 0 1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_144_531
timestamp 1
transform 1 0 49956 0 1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_144_533
timestamp 1636968456
transform 1 0 50140 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_545
timestamp 1636968456
transform 1 0 51244 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_557
timestamp 1636968456
transform 1 0 52348 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_569
timestamp 1636968456
transform 1 0 53452 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_144_581
timestamp 1
transform 1 0 54556 0 1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_144_587
timestamp 1
transform 1 0 55108 0 1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_144_589
timestamp 1636968456
transform 1 0 55292 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_601
timestamp 1636968456
transform 1 0 56396 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_613
timestamp 1636968456
transform 1 0 57500 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_625
timestamp 1636968456
transform 1 0 58604 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_144_637
timestamp 1
transform 1 0 59708 0 1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_144_643
timestamp 1
transform 1 0 60260 0 1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_144_645
timestamp 1636968456
transform 1 0 60444 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_657
timestamp 1636968456
transform 1 0 61548 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_669
timestamp 1636968456
transform 1 0 62652 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_681
timestamp 1636968456
transform 1 0 63756 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_144_693
timestamp 1
transform 1 0 64860 0 1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_144_699
timestamp 1
transform 1 0 65412 0 1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_144_701
timestamp 1636968456
transform 1 0 65596 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_713
timestamp 1636968456
transform 1 0 66700 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_725
timestamp 1636968456
transform 1 0 67804 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_737
timestamp 1636968456
transform 1 0 68908 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_144_749
timestamp 1
transform 1 0 70012 0 1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_144_755
timestamp 1
transform 1 0 70564 0 1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_144_757
timestamp 1636968456
transform 1 0 70748 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_769
timestamp 1636968456
transform 1 0 71852 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_781
timestamp 1636968456
transform 1 0 72956 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_793
timestamp 1636968456
transform 1 0 74060 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_144_805
timestamp 1
transform 1 0 75164 0 1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_144_811
timestamp 1
transform 1 0 75716 0 1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_144_813
timestamp 1636968456
transform 1 0 75900 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_825
timestamp 1636968456
transform 1 0 77004 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_837
timestamp 1636968456
transform 1 0 78108 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_849
timestamp 1636968456
transform 1 0 79212 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_144_861
timestamp 1
transform 1 0 80316 0 1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_144_867
timestamp 1
transform 1 0 80868 0 1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_144_869
timestamp 1636968456
transform 1 0 81052 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_881
timestamp 1636968456
transform 1 0 82156 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_893
timestamp 1636968456
transform 1 0 83260 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_905
timestamp 1636968456
transform 1 0 84364 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_144_917
timestamp 1
transform 1 0 85468 0 1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_144_923
timestamp 1
transform 1 0 86020 0 1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_144_925
timestamp 1636968456
transform 1 0 86204 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_937
timestamp 1636968456
transform 1 0 87308 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_949
timestamp 1636968456
transform 1 0 88412 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_961
timestamp 1636968456
transform 1 0 89516 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_144_973
timestamp 1
transform 1 0 90620 0 1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_144_979
timestamp 1
transform 1 0 91172 0 1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_144_981
timestamp 1636968456
transform 1 0 91356 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_993
timestamp 1636968456
transform 1 0 92460 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_1005
timestamp 1636968456
transform 1 0 93564 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_1017
timestamp 1636968456
transform 1 0 94668 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_144_1029
timestamp 1
transform 1 0 95772 0 1 80512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_144_1035
timestamp 1
transform 1 0 96324 0 1 80512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_144_1037
timestamp 1636968456
transform 1 0 96508 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_1049
timestamp 1636968456
transform 1 0 97612 0 1 80512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_1061
timestamp 1636968456
transform 1 0 98716 0 1 80512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_144_1073
timestamp 1
transform 1 0 99820 0 1 80512
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_145_3
timestamp 1636968456
transform 1 0 1380 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_15
timestamp 1636968456
transform 1 0 2484 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_27
timestamp 1636968456
transform 1 0 3588 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_39
timestamp 1636968456
transform 1 0 4692 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_145_51
timestamp 1
transform 1 0 5796 0 -1 81600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_145_55
timestamp 1
transform 1 0 6164 0 -1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_145_57
timestamp 1636968456
transform 1 0 6348 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_69
timestamp 1636968456
transform 1 0 7452 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_81
timestamp 1636968456
transform 1 0 8556 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_93
timestamp 1636968456
transform 1 0 9660 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_145_105
timestamp 1
transform 1 0 10764 0 -1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_145_111
timestamp 1
transform 1 0 11316 0 -1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_145_113
timestamp 1636968456
transform 1 0 11500 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_125
timestamp 1636968456
transform 1 0 12604 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_137
timestamp 1636968456
transform 1 0 13708 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_149
timestamp 1636968456
transform 1 0 14812 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_145_161
timestamp 1
transform 1 0 15916 0 -1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_145_167
timestamp 1
transform 1 0 16468 0 -1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_145_169
timestamp 1636968456
transform 1 0 16652 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_181
timestamp 1636968456
transform 1 0 17756 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_193
timestamp 1636968456
transform 1 0 18860 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_205
timestamp 1636968456
transform 1 0 19964 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_145_217
timestamp 1
transform 1 0 21068 0 -1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_145_223
timestamp 1
transform 1 0 21620 0 -1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_145_225
timestamp 1636968456
transform 1 0 21804 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_237
timestamp 1636968456
transform 1 0 22908 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_249
timestamp 1636968456
transform 1 0 24012 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_261
timestamp 1636968456
transform 1 0 25116 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_145_273
timestamp 1
transform 1 0 26220 0 -1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_145_279
timestamp 1
transform 1 0 26772 0 -1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_145_281
timestamp 1636968456
transform 1 0 26956 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_293
timestamp 1636968456
transform 1 0 28060 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_305
timestamp 1636968456
transform 1 0 29164 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_317
timestamp 1636968456
transform 1 0 30268 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_145_329
timestamp 1
transform 1 0 31372 0 -1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_145_335
timestamp 1
transform 1 0 31924 0 -1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_145_337
timestamp 1636968456
transform 1 0 32108 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_349
timestamp 1636968456
transform 1 0 33212 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_361
timestamp 1636968456
transform 1 0 34316 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_373
timestamp 1636968456
transform 1 0 35420 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_145_385
timestamp 1
transform 1 0 36524 0 -1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_145_391
timestamp 1
transform 1 0 37076 0 -1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_145_393
timestamp 1636968456
transform 1 0 37260 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_405
timestamp 1636968456
transform 1 0 38364 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_417
timestamp 1636968456
transform 1 0 39468 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_429
timestamp 1636968456
transform 1 0 40572 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_145_441
timestamp 1
transform 1 0 41676 0 -1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_145_447
timestamp 1
transform 1 0 42228 0 -1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_145_449
timestamp 1636968456
transform 1 0 42412 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_461
timestamp 1636968456
transform 1 0 43516 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_473
timestamp 1636968456
transform 1 0 44620 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_485
timestamp 1636968456
transform 1 0 45724 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_145_497
timestamp 1
transform 1 0 46828 0 -1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_145_503
timestamp 1
transform 1 0 47380 0 -1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_145_505
timestamp 1636968456
transform 1 0 47564 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_517
timestamp 1636968456
transform 1 0 48668 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_529
timestamp 1636968456
transform 1 0 49772 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_541
timestamp 1636968456
transform 1 0 50876 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_145_553
timestamp 1
transform 1 0 51980 0 -1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_145_559
timestamp 1
transform 1 0 52532 0 -1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_145_561
timestamp 1636968456
transform 1 0 52716 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_573
timestamp 1636968456
transform 1 0 53820 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_585
timestamp 1636968456
transform 1 0 54924 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_597
timestamp 1636968456
transform 1 0 56028 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_145_609
timestamp 1
transform 1 0 57132 0 -1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_145_615
timestamp 1
transform 1 0 57684 0 -1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_145_617
timestamp 1636968456
transform 1 0 57868 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_629
timestamp 1636968456
transform 1 0 58972 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_641
timestamp 1636968456
transform 1 0 60076 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_653
timestamp 1636968456
transform 1 0 61180 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_145_665
timestamp 1
transform 1 0 62284 0 -1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_145_671
timestamp 1
transform 1 0 62836 0 -1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_145_673
timestamp 1636968456
transform 1 0 63020 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_685
timestamp 1636968456
transform 1 0 64124 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_697
timestamp 1636968456
transform 1 0 65228 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_709
timestamp 1636968456
transform 1 0 66332 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_145_721
timestamp 1
transform 1 0 67436 0 -1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_145_727
timestamp 1
transform 1 0 67988 0 -1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_145_729
timestamp 1636968456
transform 1 0 68172 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_741
timestamp 1636968456
transform 1 0 69276 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_753
timestamp 1636968456
transform 1 0 70380 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_765
timestamp 1636968456
transform 1 0 71484 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_145_777
timestamp 1
transform 1 0 72588 0 -1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_145_783
timestamp 1
transform 1 0 73140 0 -1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_145_785
timestamp 1636968456
transform 1 0 73324 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_797
timestamp 1636968456
transform 1 0 74428 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_809
timestamp 1636968456
transform 1 0 75532 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_821
timestamp 1636968456
transform 1 0 76636 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_145_833
timestamp 1
transform 1 0 77740 0 -1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_145_839
timestamp 1
transform 1 0 78292 0 -1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_145_841
timestamp 1636968456
transform 1 0 78476 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_853
timestamp 1636968456
transform 1 0 79580 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_865
timestamp 1636968456
transform 1 0 80684 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_877
timestamp 1636968456
transform 1 0 81788 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_145_889
timestamp 1
transform 1 0 82892 0 -1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_145_895
timestamp 1
transform 1 0 83444 0 -1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_145_897
timestamp 1636968456
transform 1 0 83628 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_909
timestamp 1636968456
transform 1 0 84732 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_921
timestamp 1636968456
transform 1 0 85836 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_933
timestamp 1636968456
transform 1 0 86940 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_145_945
timestamp 1
transform 1 0 88044 0 -1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_145_951
timestamp 1
transform 1 0 88596 0 -1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_145_953
timestamp 1636968456
transform 1 0 88780 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_965
timestamp 1636968456
transform 1 0 89884 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_977
timestamp 1636968456
transform 1 0 90988 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_989
timestamp 1636968456
transform 1 0 92092 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_145_1001
timestamp 1
transform 1 0 93196 0 -1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_145_1007
timestamp 1
transform 1 0 93748 0 -1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_145_1009
timestamp 1636968456
transform 1 0 93932 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_1021
timestamp 1636968456
transform 1 0 95036 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_1033
timestamp 1636968456
transform 1 0 96140 0 -1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_1045
timestamp 1636968456
transform 1 0 97244 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_145_1057
timestamp 1
transform 1 0 98348 0 -1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_145_1063
timestamp 1
transform 1 0 98900 0 -1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_145_1065
timestamp 1636968456
transform 1 0 99084 0 -1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_145_1077
timestamp 1
transform 1 0 100188 0 -1 81600
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_146_3
timestamp 1636968456
transform 1 0 1380 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_15
timestamp 1636968456
transform 1 0 2484 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_146_27
timestamp 1
transform 1 0 3588 0 1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_146_29
timestamp 1636968456
transform 1 0 3772 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_41
timestamp 1636968456
transform 1 0 4876 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_53
timestamp 1636968456
transform 1 0 5980 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_65
timestamp 1636968456
transform 1 0 7084 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_146_77
timestamp 1
transform 1 0 8188 0 1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_146_83
timestamp 1
transform 1 0 8740 0 1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_146_85
timestamp 1636968456
transform 1 0 8924 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_97
timestamp 1636968456
transform 1 0 10028 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_109
timestamp 1636968456
transform 1 0 11132 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_121
timestamp 1636968456
transform 1 0 12236 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_146_133
timestamp 1
transform 1 0 13340 0 1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_146_139
timestamp 1
transform 1 0 13892 0 1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_146_141
timestamp 1636968456
transform 1 0 14076 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_153
timestamp 1636968456
transform 1 0 15180 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_165
timestamp 1636968456
transform 1 0 16284 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_177
timestamp 1636968456
transform 1 0 17388 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_146_189
timestamp 1
transform 1 0 18492 0 1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_146_195
timestamp 1
transform 1 0 19044 0 1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_146_197
timestamp 1636968456
transform 1 0 19228 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_209
timestamp 1636968456
transform 1 0 20332 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_221
timestamp 1636968456
transform 1 0 21436 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_233
timestamp 1636968456
transform 1 0 22540 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_146_245
timestamp 1
transform 1 0 23644 0 1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_146_251
timestamp 1
transform 1 0 24196 0 1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_146_253
timestamp 1636968456
transform 1 0 24380 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_265
timestamp 1636968456
transform 1 0 25484 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_277
timestamp 1636968456
transform 1 0 26588 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_289
timestamp 1636968456
transform 1 0 27692 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_146_301
timestamp 1
transform 1 0 28796 0 1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_146_307
timestamp 1
transform 1 0 29348 0 1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_146_309
timestamp 1636968456
transform 1 0 29532 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_321
timestamp 1636968456
transform 1 0 30636 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_333
timestamp 1636968456
transform 1 0 31740 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_345
timestamp 1636968456
transform 1 0 32844 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_146_357
timestamp 1
transform 1 0 33948 0 1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_146_363
timestamp 1
transform 1 0 34500 0 1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_146_365
timestamp 1636968456
transform 1 0 34684 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_377
timestamp 1636968456
transform 1 0 35788 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_389
timestamp 1636968456
transform 1 0 36892 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_401
timestamp 1636968456
transform 1 0 37996 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_146_413
timestamp 1
transform 1 0 39100 0 1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_146_419
timestamp 1
transform 1 0 39652 0 1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_146_421
timestamp 1636968456
transform 1 0 39836 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_433
timestamp 1636968456
transform 1 0 40940 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_445
timestamp 1636968456
transform 1 0 42044 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_457
timestamp 1636968456
transform 1 0 43148 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_146_469
timestamp 1
transform 1 0 44252 0 1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_146_475
timestamp 1
transform 1 0 44804 0 1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_146_477
timestamp 1636968456
transform 1 0 44988 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_489
timestamp 1636968456
transform 1 0 46092 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_501
timestamp 1636968456
transform 1 0 47196 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_513
timestamp 1636968456
transform 1 0 48300 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_146_525
timestamp 1
transform 1 0 49404 0 1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_146_531
timestamp 1
transform 1 0 49956 0 1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_146_533
timestamp 1636968456
transform 1 0 50140 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_545
timestamp 1636968456
transform 1 0 51244 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_557
timestamp 1636968456
transform 1 0 52348 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_569
timestamp 1636968456
transform 1 0 53452 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_146_581
timestamp 1
transform 1 0 54556 0 1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_146_587
timestamp 1
transform 1 0 55108 0 1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_146_589
timestamp 1636968456
transform 1 0 55292 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_601
timestamp 1636968456
transform 1 0 56396 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_613
timestamp 1636968456
transform 1 0 57500 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_625
timestamp 1636968456
transform 1 0 58604 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_146_637
timestamp 1
transform 1 0 59708 0 1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_146_643
timestamp 1
transform 1 0 60260 0 1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_146_645
timestamp 1636968456
transform 1 0 60444 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_657
timestamp 1636968456
transform 1 0 61548 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_669
timestamp 1636968456
transform 1 0 62652 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_681
timestamp 1636968456
transform 1 0 63756 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_146_693
timestamp 1
transform 1 0 64860 0 1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_146_699
timestamp 1
transform 1 0 65412 0 1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_146_701
timestamp 1636968456
transform 1 0 65596 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_713
timestamp 1636968456
transform 1 0 66700 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_725
timestamp 1636968456
transform 1 0 67804 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_737
timestamp 1636968456
transform 1 0 68908 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_146_749
timestamp 1
transform 1 0 70012 0 1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_146_755
timestamp 1
transform 1 0 70564 0 1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_146_757
timestamp 1636968456
transform 1 0 70748 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_769
timestamp 1636968456
transform 1 0 71852 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_781
timestamp 1636968456
transform 1 0 72956 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_793
timestamp 1636968456
transform 1 0 74060 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_146_805
timestamp 1
transform 1 0 75164 0 1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_146_811
timestamp 1
transform 1 0 75716 0 1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_146_813
timestamp 1636968456
transform 1 0 75900 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_825
timestamp 1636968456
transform 1 0 77004 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_837
timestamp 1636968456
transform 1 0 78108 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_849
timestamp 1636968456
transform 1 0 79212 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_146_861
timestamp 1
transform 1 0 80316 0 1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_146_867
timestamp 1
transform 1 0 80868 0 1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_146_869
timestamp 1636968456
transform 1 0 81052 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_881
timestamp 1636968456
transform 1 0 82156 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_893
timestamp 1636968456
transform 1 0 83260 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_905
timestamp 1636968456
transform 1 0 84364 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_146_917
timestamp 1
transform 1 0 85468 0 1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_146_923
timestamp 1
transform 1 0 86020 0 1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_146_925
timestamp 1636968456
transform 1 0 86204 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_937
timestamp 1636968456
transform 1 0 87308 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_949
timestamp 1636968456
transform 1 0 88412 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_961
timestamp 1636968456
transform 1 0 89516 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_146_973
timestamp 1
transform 1 0 90620 0 1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_146_979
timestamp 1
transform 1 0 91172 0 1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_146_981
timestamp 1636968456
transform 1 0 91356 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_993
timestamp 1636968456
transform 1 0 92460 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_1005
timestamp 1636968456
transform 1 0 93564 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_1017
timestamp 1636968456
transform 1 0 94668 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_146_1029
timestamp 1
transform 1 0 95772 0 1 81600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_146_1035
timestamp 1
transform 1 0 96324 0 1 81600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_146_1037
timestamp 1636968456
transform 1 0 96508 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_1049
timestamp 1636968456
transform 1 0 97612 0 1 81600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_1061
timestamp 1636968456
transform 1 0 98716 0 1 81600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_146_1073
timestamp 1
transform 1 0 99820 0 1 81600
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_147_3
timestamp 1636968456
transform 1 0 1380 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_15
timestamp 1636968456
transform 1 0 2484 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_27
timestamp 1636968456
transform 1 0 3588 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_39
timestamp 1636968456
transform 1 0 4692 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_147_51
timestamp 1
transform 1 0 5796 0 -1 82688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_147_55
timestamp 1
transform 1 0 6164 0 -1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_147_57
timestamp 1636968456
transform 1 0 6348 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_69
timestamp 1636968456
transform 1 0 7452 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_81
timestamp 1636968456
transform 1 0 8556 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_93
timestamp 1636968456
transform 1 0 9660 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_147_105
timestamp 1
transform 1 0 10764 0 -1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_147_111
timestamp 1
transform 1 0 11316 0 -1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_147_113
timestamp 1636968456
transform 1 0 11500 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_125
timestamp 1636968456
transform 1 0 12604 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_137
timestamp 1636968456
transform 1 0 13708 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_149
timestamp 1636968456
transform 1 0 14812 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_147_161
timestamp 1
transform 1 0 15916 0 -1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_147_167
timestamp 1
transform 1 0 16468 0 -1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_147_169
timestamp 1636968456
transform 1 0 16652 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_181
timestamp 1636968456
transform 1 0 17756 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_193
timestamp 1636968456
transform 1 0 18860 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_205
timestamp 1636968456
transform 1 0 19964 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_147_217
timestamp 1
transform 1 0 21068 0 -1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_147_223
timestamp 1
transform 1 0 21620 0 -1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_147_225
timestamp 1636968456
transform 1 0 21804 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_237
timestamp 1636968456
transform 1 0 22908 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_249
timestamp 1636968456
transform 1 0 24012 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_261
timestamp 1636968456
transform 1 0 25116 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_147_273
timestamp 1
transform 1 0 26220 0 -1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_147_279
timestamp 1
transform 1 0 26772 0 -1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_147_281
timestamp 1636968456
transform 1 0 26956 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_293
timestamp 1636968456
transform 1 0 28060 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_305
timestamp 1636968456
transform 1 0 29164 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_317
timestamp 1636968456
transform 1 0 30268 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_147_329
timestamp 1
transform 1 0 31372 0 -1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_147_335
timestamp 1
transform 1 0 31924 0 -1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_147_337
timestamp 1636968456
transform 1 0 32108 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_349
timestamp 1636968456
transform 1 0 33212 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_361
timestamp 1636968456
transform 1 0 34316 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_373
timestamp 1636968456
transform 1 0 35420 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_147_385
timestamp 1
transform 1 0 36524 0 -1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_147_391
timestamp 1
transform 1 0 37076 0 -1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_147_393
timestamp 1636968456
transform 1 0 37260 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_405
timestamp 1636968456
transform 1 0 38364 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_417
timestamp 1636968456
transform 1 0 39468 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_429
timestamp 1636968456
transform 1 0 40572 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_147_441
timestamp 1
transform 1 0 41676 0 -1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_147_447
timestamp 1
transform 1 0 42228 0 -1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_147_449
timestamp 1636968456
transform 1 0 42412 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_461
timestamp 1636968456
transform 1 0 43516 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_473
timestamp 1636968456
transform 1 0 44620 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_485
timestamp 1636968456
transform 1 0 45724 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_147_497
timestamp 1
transform 1 0 46828 0 -1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_147_503
timestamp 1
transform 1 0 47380 0 -1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_147_505
timestamp 1636968456
transform 1 0 47564 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_517
timestamp 1636968456
transform 1 0 48668 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_529
timestamp 1636968456
transform 1 0 49772 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_541
timestamp 1636968456
transform 1 0 50876 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_147_553
timestamp 1
transform 1 0 51980 0 -1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_147_559
timestamp 1
transform 1 0 52532 0 -1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_147_561
timestamp 1636968456
transform 1 0 52716 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_573
timestamp 1636968456
transform 1 0 53820 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_585
timestamp 1636968456
transform 1 0 54924 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_597
timestamp 1636968456
transform 1 0 56028 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_147_609
timestamp 1
transform 1 0 57132 0 -1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_147_615
timestamp 1
transform 1 0 57684 0 -1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_147_617
timestamp 1636968456
transform 1 0 57868 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_629
timestamp 1636968456
transform 1 0 58972 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_641
timestamp 1636968456
transform 1 0 60076 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_653
timestamp 1636968456
transform 1 0 61180 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_147_665
timestamp 1
transform 1 0 62284 0 -1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_147_671
timestamp 1
transform 1 0 62836 0 -1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_147_673
timestamp 1636968456
transform 1 0 63020 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_685
timestamp 1636968456
transform 1 0 64124 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_697
timestamp 1636968456
transform 1 0 65228 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_709
timestamp 1636968456
transform 1 0 66332 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_147_721
timestamp 1
transform 1 0 67436 0 -1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_147_727
timestamp 1
transform 1 0 67988 0 -1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_147_729
timestamp 1636968456
transform 1 0 68172 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_741
timestamp 1636968456
transform 1 0 69276 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_753
timestamp 1636968456
transform 1 0 70380 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_765
timestamp 1636968456
transform 1 0 71484 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_147_777
timestamp 1
transform 1 0 72588 0 -1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_147_783
timestamp 1
transform 1 0 73140 0 -1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_147_785
timestamp 1636968456
transform 1 0 73324 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_797
timestamp 1636968456
transform 1 0 74428 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_809
timestamp 1636968456
transform 1 0 75532 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_821
timestamp 1636968456
transform 1 0 76636 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_147_833
timestamp 1
transform 1 0 77740 0 -1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_147_839
timestamp 1
transform 1 0 78292 0 -1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_147_841
timestamp 1636968456
transform 1 0 78476 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_853
timestamp 1636968456
transform 1 0 79580 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_865
timestamp 1636968456
transform 1 0 80684 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_877
timestamp 1636968456
transform 1 0 81788 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_147_889
timestamp 1
transform 1 0 82892 0 -1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_147_895
timestamp 1
transform 1 0 83444 0 -1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_147_897
timestamp 1636968456
transform 1 0 83628 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_909
timestamp 1636968456
transform 1 0 84732 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_921
timestamp 1636968456
transform 1 0 85836 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_933
timestamp 1636968456
transform 1 0 86940 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_147_945
timestamp 1
transform 1 0 88044 0 -1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_147_951
timestamp 1
transform 1 0 88596 0 -1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_147_953
timestamp 1636968456
transform 1 0 88780 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_965
timestamp 1636968456
transform 1 0 89884 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_977
timestamp 1636968456
transform 1 0 90988 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_989
timestamp 1636968456
transform 1 0 92092 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_147_1001
timestamp 1
transform 1 0 93196 0 -1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_147_1007
timestamp 1
transform 1 0 93748 0 -1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_147_1009
timestamp 1636968456
transform 1 0 93932 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_1021
timestamp 1636968456
transform 1 0 95036 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_1033
timestamp 1636968456
transform 1 0 96140 0 -1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_1045
timestamp 1636968456
transform 1 0 97244 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_147_1057
timestamp 1
transform 1 0 98348 0 -1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_147_1063
timestamp 1
transform 1 0 98900 0 -1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_147_1065
timestamp 1636968456
transform 1 0 99084 0 -1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_147_1077
timestamp 1
transform 1 0 100188 0 -1 82688
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_148_3
timestamp 1636968456
transform 1 0 1380 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_15
timestamp 1636968456
transform 1 0 2484 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_148_27
timestamp 1
transform 1 0 3588 0 1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_148_29
timestamp 1636968456
transform 1 0 3772 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_41
timestamp 1636968456
transform 1 0 4876 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_53
timestamp 1636968456
transform 1 0 5980 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_65
timestamp 1636968456
transform 1 0 7084 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_148_77
timestamp 1
transform 1 0 8188 0 1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_148_83
timestamp 1
transform 1 0 8740 0 1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_148_85
timestamp 1636968456
transform 1 0 8924 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_97
timestamp 1636968456
transform 1 0 10028 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_109
timestamp 1636968456
transform 1 0 11132 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_121
timestamp 1636968456
transform 1 0 12236 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_148_133
timestamp 1
transform 1 0 13340 0 1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_148_139
timestamp 1
transform 1 0 13892 0 1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_148_141
timestamp 1636968456
transform 1 0 14076 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_153
timestamp 1636968456
transform 1 0 15180 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_165
timestamp 1636968456
transform 1 0 16284 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_177
timestamp 1636968456
transform 1 0 17388 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_148_189
timestamp 1
transform 1 0 18492 0 1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_148_195
timestamp 1
transform 1 0 19044 0 1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_148_197
timestamp 1636968456
transform 1 0 19228 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_209
timestamp 1636968456
transform 1 0 20332 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_221
timestamp 1636968456
transform 1 0 21436 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_233
timestamp 1636968456
transform 1 0 22540 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_148_245
timestamp 1
transform 1 0 23644 0 1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_148_251
timestamp 1
transform 1 0 24196 0 1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_148_253
timestamp 1636968456
transform 1 0 24380 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_265
timestamp 1636968456
transform 1 0 25484 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_277
timestamp 1636968456
transform 1 0 26588 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_289
timestamp 1636968456
transform 1 0 27692 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_148_301
timestamp 1
transform 1 0 28796 0 1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_148_307
timestamp 1
transform 1 0 29348 0 1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_148_309
timestamp 1636968456
transform 1 0 29532 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_321
timestamp 1636968456
transform 1 0 30636 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_333
timestamp 1636968456
transform 1 0 31740 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_345
timestamp 1636968456
transform 1 0 32844 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_148_357
timestamp 1
transform 1 0 33948 0 1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_148_363
timestamp 1
transform 1 0 34500 0 1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_148_365
timestamp 1636968456
transform 1 0 34684 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_377
timestamp 1636968456
transform 1 0 35788 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_389
timestamp 1636968456
transform 1 0 36892 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_401
timestamp 1636968456
transform 1 0 37996 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_148_413
timestamp 1
transform 1 0 39100 0 1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_148_419
timestamp 1
transform 1 0 39652 0 1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_148_421
timestamp 1636968456
transform 1 0 39836 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_433
timestamp 1636968456
transform 1 0 40940 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_445
timestamp 1636968456
transform 1 0 42044 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_457
timestamp 1636968456
transform 1 0 43148 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_148_469
timestamp 1
transform 1 0 44252 0 1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_148_475
timestamp 1
transform 1 0 44804 0 1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_148_477
timestamp 1636968456
transform 1 0 44988 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_489
timestamp 1636968456
transform 1 0 46092 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_501
timestamp 1636968456
transform 1 0 47196 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_513
timestamp 1636968456
transform 1 0 48300 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_148_525
timestamp 1
transform 1 0 49404 0 1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_148_531
timestamp 1
transform 1 0 49956 0 1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_148_533
timestamp 1636968456
transform 1 0 50140 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_545
timestamp 1636968456
transform 1 0 51244 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_557
timestamp 1636968456
transform 1 0 52348 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_569
timestamp 1636968456
transform 1 0 53452 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_148_581
timestamp 1
transform 1 0 54556 0 1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_148_587
timestamp 1
transform 1 0 55108 0 1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_148_589
timestamp 1636968456
transform 1 0 55292 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_601
timestamp 1636968456
transform 1 0 56396 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_613
timestamp 1636968456
transform 1 0 57500 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_625
timestamp 1636968456
transform 1 0 58604 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_148_637
timestamp 1
transform 1 0 59708 0 1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_148_643
timestamp 1
transform 1 0 60260 0 1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_148_645
timestamp 1636968456
transform 1 0 60444 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_657
timestamp 1636968456
transform 1 0 61548 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_669
timestamp 1636968456
transform 1 0 62652 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_681
timestamp 1636968456
transform 1 0 63756 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_148_693
timestamp 1
transform 1 0 64860 0 1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_148_699
timestamp 1
transform 1 0 65412 0 1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_148_701
timestamp 1636968456
transform 1 0 65596 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_713
timestamp 1636968456
transform 1 0 66700 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_725
timestamp 1636968456
transform 1 0 67804 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_737
timestamp 1636968456
transform 1 0 68908 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_148_749
timestamp 1
transform 1 0 70012 0 1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_148_755
timestamp 1
transform 1 0 70564 0 1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_148_757
timestamp 1636968456
transform 1 0 70748 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_769
timestamp 1636968456
transform 1 0 71852 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_781
timestamp 1636968456
transform 1 0 72956 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_793
timestamp 1636968456
transform 1 0 74060 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_148_805
timestamp 1
transform 1 0 75164 0 1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_148_811
timestamp 1
transform 1 0 75716 0 1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_148_813
timestamp 1636968456
transform 1 0 75900 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_825
timestamp 1636968456
transform 1 0 77004 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_837
timestamp 1636968456
transform 1 0 78108 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_849
timestamp 1636968456
transform 1 0 79212 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_148_861
timestamp 1
transform 1 0 80316 0 1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_148_867
timestamp 1
transform 1 0 80868 0 1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_148_869
timestamp 1636968456
transform 1 0 81052 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_881
timestamp 1636968456
transform 1 0 82156 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_893
timestamp 1636968456
transform 1 0 83260 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_905
timestamp 1636968456
transform 1 0 84364 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_148_917
timestamp 1
transform 1 0 85468 0 1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_148_923
timestamp 1
transform 1 0 86020 0 1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_148_925
timestamp 1636968456
transform 1 0 86204 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_937
timestamp 1636968456
transform 1 0 87308 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_949
timestamp 1636968456
transform 1 0 88412 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_961
timestamp 1636968456
transform 1 0 89516 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_148_973
timestamp 1
transform 1 0 90620 0 1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_148_979
timestamp 1
transform 1 0 91172 0 1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_148_981
timestamp 1636968456
transform 1 0 91356 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_993
timestamp 1636968456
transform 1 0 92460 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_1005
timestamp 1636968456
transform 1 0 93564 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_1017
timestamp 1636968456
transform 1 0 94668 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_148_1029
timestamp 1
transform 1 0 95772 0 1 82688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_148_1035
timestamp 1
transform 1 0 96324 0 1 82688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_148_1037
timestamp 1636968456
transform 1 0 96508 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_1049
timestamp 1636968456
transform 1 0 97612 0 1 82688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_1061
timestamp 1636968456
transform 1 0 98716 0 1 82688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_148_1073
timestamp 1
transform 1 0 99820 0 1 82688
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_149_3
timestamp 1636968456
transform 1 0 1380 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_15
timestamp 1636968456
transform 1 0 2484 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_27
timestamp 1636968456
transform 1 0 3588 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_39
timestamp 1636968456
transform 1 0 4692 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_149_51
timestamp 1
transform 1 0 5796 0 -1 83776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_149_55
timestamp 1
transform 1 0 6164 0 -1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_149_57
timestamp 1636968456
transform 1 0 6348 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_69
timestamp 1636968456
transform 1 0 7452 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_81
timestamp 1636968456
transform 1 0 8556 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_93
timestamp 1636968456
transform 1 0 9660 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_149_105
timestamp 1
transform 1 0 10764 0 -1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_149_111
timestamp 1
transform 1 0 11316 0 -1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_149_113
timestamp 1636968456
transform 1 0 11500 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_125
timestamp 1636968456
transform 1 0 12604 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_137
timestamp 1636968456
transform 1 0 13708 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_149
timestamp 1636968456
transform 1 0 14812 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_149_161
timestamp 1
transform 1 0 15916 0 -1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_149_167
timestamp 1
transform 1 0 16468 0 -1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_149_169
timestamp 1636968456
transform 1 0 16652 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_181
timestamp 1636968456
transform 1 0 17756 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_193
timestamp 1636968456
transform 1 0 18860 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_205
timestamp 1636968456
transform 1 0 19964 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_149_217
timestamp 1
transform 1 0 21068 0 -1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_149_223
timestamp 1
transform 1 0 21620 0 -1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_149_225
timestamp 1636968456
transform 1 0 21804 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_237
timestamp 1636968456
transform 1 0 22908 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_249
timestamp 1636968456
transform 1 0 24012 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_261
timestamp 1636968456
transform 1 0 25116 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_149_273
timestamp 1
transform 1 0 26220 0 -1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_149_279
timestamp 1
transform 1 0 26772 0 -1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_149_281
timestamp 1636968456
transform 1 0 26956 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_293
timestamp 1636968456
transform 1 0 28060 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_305
timestamp 1636968456
transform 1 0 29164 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_317
timestamp 1636968456
transform 1 0 30268 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_149_329
timestamp 1
transform 1 0 31372 0 -1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_149_335
timestamp 1
transform 1 0 31924 0 -1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_149_337
timestamp 1636968456
transform 1 0 32108 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_349
timestamp 1636968456
transform 1 0 33212 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_361
timestamp 1636968456
transform 1 0 34316 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_373
timestamp 1636968456
transform 1 0 35420 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_149_385
timestamp 1
transform 1 0 36524 0 -1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_149_391
timestamp 1
transform 1 0 37076 0 -1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_149_393
timestamp 1636968456
transform 1 0 37260 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_405
timestamp 1636968456
transform 1 0 38364 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_417
timestamp 1636968456
transform 1 0 39468 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_429
timestamp 1636968456
transform 1 0 40572 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_149_441
timestamp 1
transform 1 0 41676 0 -1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_149_447
timestamp 1
transform 1 0 42228 0 -1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_149_449
timestamp 1636968456
transform 1 0 42412 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_461
timestamp 1636968456
transform 1 0 43516 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_473
timestamp 1636968456
transform 1 0 44620 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_485
timestamp 1636968456
transform 1 0 45724 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_149_497
timestamp 1
transform 1 0 46828 0 -1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_149_503
timestamp 1
transform 1 0 47380 0 -1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_149_505
timestamp 1636968456
transform 1 0 47564 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_517
timestamp 1636968456
transform 1 0 48668 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_529
timestamp 1636968456
transform 1 0 49772 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_541
timestamp 1636968456
transform 1 0 50876 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_149_553
timestamp 1
transform 1 0 51980 0 -1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_149_559
timestamp 1
transform 1 0 52532 0 -1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_149_561
timestamp 1636968456
transform 1 0 52716 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_573
timestamp 1636968456
transform 1 0 53820 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_585
timestamp 1636968456
transform 1 0 54924 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_597
timestamp 1636968456
transform 1 0 56028 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_149_609
timestamp 1
transform 1 0 57132 0 -1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_149_615
timestamp 1
transform 1 0 57684 0 -1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_149_617
timestamp 1636968456
transform 1 0 57868 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_629
timestamp 1636968456
transform 1 0 58972 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_641
timestamp 1636968456
transform 1 0 60076 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_653
timestamp 1636968456
transform 1 0 61180 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_149_665
timestamp 1
transform 1 0 62284 0 -1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_149_671
timestamp 1
transform 1 0 62836 0 -1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_149_673
timestamp 1636968456
transform 1 0 63020 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_685
timestamp 1636968456
transform 1 0 64124 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_697
timestamp 1636968456
transform 1 0 65228 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_709
timestamp 1636968456
transform 1 0 66332 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_149_721
timestamp 1
transform 1 0 67436 0 -1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_149_727
timestamp 1
transform 1 0 67988 0 -1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_149_729
timestamp 1636968456
transform 1 0 68172 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_741
timestamp 1636968456
transform 1 0 69276 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_753
timestamp 1636968456
transform 1 0 70380 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_765
timestamp 1636968456
transform 1 0 71484 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_149_777
timestamp 1
transform 1 0 72588 0 -1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_149_783
timestamp 1
transform 1 0 73140 0 -1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_149_785
timestamp 1636968456
transform 1 0 73324 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_797
timestamp 1636968456
transform 1 0 74428 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_809
timestamp 1636968456
transform 1 0 75532 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_821
timestamp 1636968456
transform 1 0 76636 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_149_833
timestamp 1
transform 1 0 77740 0 -1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_149_839
timestamp 1
transform 1 0 78292 0 -1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_149_841
timestamp 1636968456
transform 1 0 78476 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_853
timestamp 1636968456
transform 1 0 79580 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_865
timestamp 1636968456
transform 1 0 80684 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_877
timestamp 1636968456
transform 1 0 81788 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_149_889
timestamp 1
transform 1 0 82892 0 -1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_149_895
timestamp 1
transform 1 0 83444 0 -1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_149_897
timestamp 1636968456
transform 1 0 83628 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_909
timestamp 1636968456
transform 1 0 84732 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_921
timestamp 1636968456
transform 1 0 85836 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_933
timestamp 1636968456
transform 1 0 86940 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_149_945
timestamp 1
transform 1 0 88044 0 -1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_149_951
timestamp 1
transform 1 0 88596 0 -1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_149_953
timestamp 1636968456
transform 1 0 88780 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_965
timestamp 1636968456
transform 1 0 89884 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_977
timestamp 1636968456
transform 1 0 90988 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_989
timestamp 1636968456
transform 1 0 92092 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_149_1001
timestamp 1
transform 1 0 93196 0 -1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_149_1007
timestamp 1
transform 1 0 93748 0 -1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_149_1009
timestamp 1636968456
transform 1 0 93932 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_1021
timestamp 1636968456
transform 1 0 95036 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_1033
timestamp 1636968456
transform 1 0 96140 0 -1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_1045
timestamp 1636968456
transform 1 0 97244 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_149_1057
timestamp 1
transform 1 0 98348 0 -1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_149_1063
timestamp 1
transform 1 0 98900 0 -1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_149_1065
timestamp 1636968456
transform 1 0 99084 0 -1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_149_1077
timestamp 1
transform 1 0 100188 0 -1 83776
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_150_3
timestamp 1636968456
transform 1 0 1380 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_15
timestamp 1636968456
transform 1 0 2484 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_150_27
timestamp 1
transform 1 0 3588 0 1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_150_29
timestamp 1636968456
transform 1 0 3772 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_41
timestamp 1636968456
transform 1 0 4876 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_53
timestamp 1636968456
transform 1 0 5980 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_65
timestamp 1636968456
transform 1 0 7084 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_150_77
timestamp 1
transform 1 0 8188 0 1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_150_83
timestamp 1
transform 1 0 8740 0 1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_150_85
timestamp 1636968456
transform 1 0 8924 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_97
timestamp 1636968456
transform 1 0 10028 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_109
timestamp 1636968456
transform 1 0 11132 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_121
timestamp 1636968456
transform 1 0 12236 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_150_133
timestamp 1
transform 1 0 13340 0 1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_150_139
timestamp 1
transform 1 0 13892 0 1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_150_141
timestamp 1636968456
transform 1 0 14076 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_153
timestamp 1636968456
transform 1 0 15180 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_165
timestamp 1636968456
transform 1 0 16284 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_177
timestamp 1636968456
transform 1 0 17388 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_150_189
timestamp 1
transform 1 0 18492 0 1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_150_195
timestamp 1
transform 1 0 19044 0 1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_150_197
timestamp 1636968456
transform 1 0 19228 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_209
timestamp 1636968456
transform 1 0 20332 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_221
timestamp 1636968456
transform 1 0 21436 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_233
timestamp 1636968456
transform 1 0 22540 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_150_245
timestamp 1
transform 1 0 23644 0 1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_150_251
timestamp 1
transform 1 0 24196 0 1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_150_253
timestamp 1636968456
transform 1 0 24380 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_265
timestamp 1636968456
transform 1 0 25484 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_277
timestamp 1636968456
transform 1 0 26588 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_289
timestamp 1636968456
transform 1 0 27692 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_150_301
timestamp 1
transform 1 0 28796 0 1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_150_307
timestamp 1
transform 1 0 29348 0 1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_150_309
timestamp 1636968456
transform 1 0 29532 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_321
timestamp 1636968456
transform 1 0 30636 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_333
timestamp 1636968456
transform 1 0 31740 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_345
timestamp 1636968456
transform 1 0 32844 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_150_357
timestamp 1
transform 1 0 33948 0 1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_150_363
timestamp 1
transform 1 0 34500 0 1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_150_365
timestamp 1636968456
transform 1 0 34684 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_377
timestamp 1636968456
transform 1 0 35788 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_389
timestamp 1636968456
transform 1 0 36892 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_401
timestamp 1636968456
transform 1 0 37996 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_150_413
timestamp 1
transform 1 0 39100 0 1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_150_419
timestamp 1
transform 1 0 39652 0 1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_150_421
timestamp 1636968456
transform 1 0 39836 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_433
timestamp 1636968456
transform 1 0 40940 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_445
timestamp 1636968456
transform 1 0 42044 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_457
timestamp 1636968456
transform 1 0 43148 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_150_469
timestamp 1
transform 1 0 44252 0 1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_150_475
timestamp 1
transform 1 0 44804 0 1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_150_477
timestamp 1636968456
transform 1 0 44988 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_489
timestamp 1636968456
transform 1 0 46092 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_501
timestamp 1636968456
transform 1 0 47196 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_513
timestamp 1636968456
transform 1 0 48300 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_150_525
timestamp 1
transform 1 0 49404 0 1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_150_531
timestamp 1
transform 1 0 49956 0 1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_150_533
timestamp 1636968456
transform 1 0 50140 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_545
timestamp 1636968456
transform 1 0 51244 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_557
timestamp 1636968456
transform 1 0 52348 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_569
timestamp 1636968456
transform 1 0 53452 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_150_581
timestamp 1
transform 1 0 54556 0 1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_150_587
timestamp 1
transform 1 0 55108 0 1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_150_589
timestamp 1636968456
transform 1 0 55292 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_601
timestamp 1636968456
transform 1 0 56396 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_613
timestamp 1636968456
transform 1 0 57500 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_625
timestamp 1636968456
transform 1 0 58604 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_150_637
timestamp 1
transform 1 0 59708 0 1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_150_643
timestamp 1
transform 1 0 60260 0 1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_150_645
timestamp 1636968456
transform 1 0 60444 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_657
timestamp 1636968456
transform 1 0 61548 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_669
timestamp 1636968456
transform 1 0 62652 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_681
timestamp 1636968456
transform 1 0 63756 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_150_693
timestamp 1
transform 1 0 64860 0 1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_150_699
timestamp 1
transform 1 0 65412 0 1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_150_701
timestamp 1636968456
transform 1 0 65596 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_713
timestamp 1636968456
transform 1 0 66700 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_725
timestamp 1636968456
transform 1 0 67804 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_737
timestamp 1636968456
transform 1 0 68908 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_150_749
timestamp 1
transform 1 0 70012 0 1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_150_755
timestamp 1
transform 1 0 70564 0 1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_150_757
timestamp 1636968456
transform 1 0 70748 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_769
timestamp 1636968456
transform 1 0 71852 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_781
timestamp 1636968456
transform 1 0 72956 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_793
timestamp 1636968456
transform 1 0 74060 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_150_805
timestamp 1
transform 1 0 75164 0 1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_150_811
timestamp 1
transform 1 0 75716 0 1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_150_813
timestamp 1636968456
transform 1 0 75900 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_825
timestamp 1636968456
transform 1 0 77004 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_837
timestamp 1636968456
transform 1 0 78108 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_849
timestamp 1636968456
transform 1 0 79212 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_150_861
timestamp 1
transform 1 0 80316 0 1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_150_867
timestamp 1
transform 1 0 80868 0 1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_150_869
timestamp 1636968456
transform 1 0 81052 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_881
timestamp 1636968456
transform 1 0 82156 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_893
timestamp 1636968456
transform 1 0 83260 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_905
timestamp 1636968456
transform 1 0 84364 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_150_917
timestamp 1
transform 1 0 85468 0 1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_150_923
timestamp 1
transform 1 0 86020 0 1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_150_925
timestamp 1636968456
transform 1 0 86204 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_937
timestamp 1636968456
transform 1 0 87308 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_949
timestamp 1636968456
transform 1 0 88412 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_961
timestamp 1636968456
transform 1 0 89516 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_150_973
timestamp 1
transform 1 0 90620 0 1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_150_979
timestamp 1
transform 1 0 91172 0 1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_150_981
timestamp 1636968456
transform 1 0 91356 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_993
timestamp 1636968456
transform 1 0 92460 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_1005
timestamp 1636968456
transform 1 0 93564 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_1017
timestamp 1636968456
transform 1 0 94668 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_150_1029
timestamp 1
transform 1 0 95772 0 1 83776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_150_1035
timestamp 1
transform 1 0 96324 0 1 83776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_150_1037
timestamp 1636968456
transform 1 0 96508 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_1049
timestamp 1636968456
transform 1 0 97612 0 1 83776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_1061
timestamp 1636968456
transform 1 0 98716 0 1 83776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_150_1073
timestamp 1
transform 1 0 99820 0 1 83776
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_151_3
timestamp 1636968456
transform 1 0 1380 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_15
timestamp 1636968456
transform 1 0 2484 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_27
timestamp 1636968456
transform 1 0 3588 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_39
timestamp 1636968456
transform 1 0 4692 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_151_51
timestamp 1
transform 1 0 5796 0 -1 84864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_151_55
timestamp 1
transform 1 0 6164 0 -1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_151_57
timestamp 1636968456
transform 1 0 6348 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_69
timestamp 1636968456
transform 1 0 7452 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_81
timestamp 1636968456
transform 1 0 8556 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_93
timestamp 1636968456
transform 1 0 9660 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_151_105
timestamp 1
transform 1 0 10764 0 -1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_151_111
timestamp 1
transform 1 0 11316 0 -1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_151_113
timestamp 1636968456
transform 1 0 11500 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_125
timestamp 1636968456
transform 1 0 12604 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_137
timestamp 1636968456
transform 1 0 13708 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_149
timestamp 1636968456
transform 1 0 14812 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_151_161
timestamp 1
transform 1 0 15916 0 -1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_151_167
timestamp 1
transform 1 0 16468 0 -1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_151_169
timestamp 1636968456
transform 1 0 16652 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_181
timestamp 1636968456
transform 1 0 17756 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_193
timestamp 1636968456
transform 1 0 18860 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_205
timestamp 1636968456
transform 1 0 19964 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_151_217
timestamp 1
transform 1 0 21068 0 -1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_151_223
timestamp 1
transform 1 0 21620 0 -1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_151_225
timestamp 1636968456
transform 1 0 21804 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_237
timestamp 1636968456
transform 1 0 22908 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_249
timestamp 1636968456
transform 1 0 24012 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_261
timestamp 1636968456
transform 1 0 25116 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_151_273
timestamp 1
transform 1 0 26220 0 -1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_151_279
timestamp 1
transform 1 0 26772 0 -1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_151_281
timestamp 1636968456
transform 1 0 26956 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_293
timestamp 1636968456
transform 1 0 28060 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_305
timestamp 1636968456
transform 1 0 29164 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_317
timestamp 1636968456
transform 1 0 30268 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_151_329
timestamp 1
transform 1 0 31372 0 -1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_151_335
timestamp 1
transform 1 0 31924 0 -1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_151_337
timestamp 1636968456
transform 1 0 32108 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_349
timestamp 1636968456
transform 1 0 33212 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_361
timestamp 1636968456
transform 1 0 34316 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_373
timestamp 1636968456
transform 1 0 35420 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_151_385
timestamp 1
transform 1 0 36524 0 -1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_151_391
timestamp 1
transform 1 0 37076 0 -1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_151_393
timestamp 1636968456
transform 1 0 37260 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_405
timestamp 1636968456
transform 1 0 38364 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_417
timestamp 1636968456
transform 1 0 39468 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_429
timestamp 1636968456
transform 1 0 40572 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_151_441
timestamp 1
transform 1 0 41676 0 -1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_151_447
timestamp 1
transform 1 0 42228 0 -1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_151_449
timestamp 1636968456
transform 1 0 42412 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_461
timestamp 1636968456
transform 1 0 43516 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_473
timestamp 1636968456
transform 1 0 44620 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_485
timestamp 1636968456
transform 1 0 45724 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_151_497
timestamp 1
transform 1 0 46828 0 -1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_151_503
timestamp 1
transform 1 0 47380 0 -1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_151_505
timestamp 1636968456
transform 1 0 47564 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_517
timestamp 1636968456
transform 1 0 48668 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_529
timestamp 1636968456
transform 1 0 49772 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_541
timestamp 1636968456
transform 1 0 50876 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_151_553
timestamp 1
transform 1 0 51980 0 -1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_151_559
timestamp 1
transform 1 0 52532 0 -1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_151_561
timestamp 1636968456
transform 1 0 52716 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_573
timestamp 1636968456
transform 1 0 53820 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_585
timestamp 1636968456
transform 1 0 54924 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_597
timestamp 1636968456
transform 1 0 56028 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_151_609
timestamp 1
transform 1 0 57132 0 -1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_151_615
timestamp 1
transform 1 0 57684 0 -1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_151_617
timestamp 1636968456
transform 1 0 57868 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_629
timestamp 1636968456
transform 1 0 58972 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_641
timestamp 1636968456
transform 1 0 60076 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_653
timestamp 1636968456
transform 1 0 61180 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_151_665
timestamp 1
transform 1 0 62284 0 -1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_151_671
timestamp 1
transform 1 0 62836 0 -1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_151_673
timestamp 1636968456
transform 1 0 63020 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_685
timestamp 1636968456
transform 1 0 64124 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_697
timestamp 1636968456
transform 1 0 65228 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_709
timestamp 1636968456
transform 1 0 66332 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_151_721
timestamp 1
transform 1 0 67436 0 -1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_151_727
timestamp 1
transform 1 0 67988 0 -1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_151_729
timestamp 1636968456
transform 1 0 68172 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_741
timestamp 1636968456
transform 1 0 69276 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_753
timestamp 1636968456
transform 1 0 70380 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_765
timestamp 1636968456
transform 1 0 71484 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_151_777
timestamp 1
transform 1 0 72588 0 -1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_151_783
timestamp 1
transform 1 0 73140 0 -1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_151_785
timestamp 1636968456
transform 1 0 73324 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_797
timestamp 1636968456
transform 1 0 74428 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_809
timestamp 1636968456
transform 1 0 75532 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_821
timestamp 1636968456
transform 1 0 76636 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_151_833
timestamp 1
transform 1 0 77740 0 -1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_151_839
timestamp 1
transform 1 0 78292 0 -1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_151_841
timestamp 1636968456
transform 1 0 78476 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_853
timestamp 1636968456
transform 1 0 79580 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_865
timestamp 1636968456
transform 1 0 80684 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_877
timestamp 1636968456
transform 1 0 81788 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_151_889
timestamp 1
transform 1 0 82892 0 -1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_151_895
timestamp 1
transform 1 0 83444 0 -1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_151_897
timestamp 1636968456
transform 1 0 83628 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_909
timestamp 1636968456
transform 1 0 84732 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_921
timestamp 1636968456
transform 1 0 85836 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_933
timestamp 1636968456
transform 1 0 86940 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_151_945
timestamp 1
transform 1 0 88044 0 -1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_151_951
timestamp 1
transform 1 0 88596 0 -1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_151_953
timestamp 1636968456
transform 1 0 88780 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_965
timestamp 1636968456
transform 1 0 89884 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_977
timestamp 1636968456
transform 1 0 90988 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_989
timestamp 1636968456
transform 1 0 92092 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_151_1001
timestamp 1
transform 1 0 93196 0 -1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_151_1007
timestamp 1
transform 1 0 93748 0 -1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_151_1009
timestamp 1636968456
transform 1 0 93932 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_1021
timestamp 1636968456
transform 1 0 95036 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_1033
timestamp 1636968456
transform 1 0 96140 0 -1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_1045
timestamp 1636968456
transform 1 0 97244 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_151_1057
timestamp 1
transform 1 0 98348 0 -1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_151_1063
timestamp 1
transform 1 0 98900 0 -1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_151_1065
timestamp 1636968456
transform 1 0 99084 0 -1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_151_1077
timestamp 1
transform 1 0 100188 0 -1 84864
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_152_3
timestamp 1636968456
transform 1 0 1380 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_15
timestamp 1636968456
transform 1 0 2484 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_152_27
timestamp 1
transform 1 0 3588 0 1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_152_29
timestamp 1636968456
transform 1 0 3772 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_41
timestamp 1636968456
transform 1 0 4876 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_53
timestamp 1636968456
transform 1 0 5980 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_65
timestamp 1636968456
transform 1 0 7084 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_152_77
timestamp 1
transform 1 0 8188 0 1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_152_83
timestamp 1
transform 1 0 8740 0 1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_152_85
timestamp 1636968456
transform 1 0 8924 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_97
timestamp 1636968456
transform 1 0 10028 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_109
timestamp 1636968456
transform 1 0 11132 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_121
timestamp 1636968456
transform 1 0 12236 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_152_133
timestamp 1
transform 1 0 13340 0 1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_152_139
timestamp 1
transform 1 0 13892 0 1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_152_141
timestamp 1636968456
transform 1 0 14076 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_153
timestamp 1636968456
transform 1 0 15180 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_165
timestamp 1636968456
transform 1 0 16284 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_177
timestamp 1636968456
transform 1 0 17388 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_152_189
timestamp 1
transform 1 0 18492 0 1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_152_195
timestamp 1
transform 1 0 19044 0 1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_152_197
timestamp 1636968456
transform 1 0 19228 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_209
timestamp 1636968456
transform 1 0 20332 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_221
timestamp 1636968456
transform 1 0 21436 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_233
timestamp 1636968456
transform 1 0 22540 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_152_245
timestamp 1
transform 1 0 23644 0 1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_152_251
timestamp 1
transform 1 0 24196 0 1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_152_253
timestamp 1636968456
transform 1 0 24380 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_265
timestamp 1636968456
transform 1 0 25484 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_277
timestamp 1636968456
transform 1 0 26588 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_289
timestamp 1636968456
transform 1 0 27692 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_152_301
timestamp 1
transform 1 0 28796 0 1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_152_307
timestamp 1
transform 1 0 29348 0 1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_152_309
timestamp 1636968456
transform 1 0 29532 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_321
timestamp 1636968456
transform 1 0 30636 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_333
timestamp 1636968456
transform 1 0 31740 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_345
timestamp 1636968456
transform 1 0 32844 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_152_357
timestamp 1
transform 1 0 33948 0 1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_152_363
timestamp 1
transform 1 0 34500 0 1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_152_365
timestamp 1636968456
transform 1 0 34684 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_377
timestamp 1636968456
transform 1 0 35788 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_389
timestamp 1636968456
transform 1 0 36892 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_401
timestamp 1636968456
transform 1 0 37996 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_152_413
timestamp 1
transform 1 0 39100 0 1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_152_419
timestamp 1
transform 1 0 39652 0 1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_152_421
timestamp 1636968456
transform 1 0 39836 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_433
timestamp 1636968456
transform 1 0 40940 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_445
timestamp 1636968456
transform 1 0 42044 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_457
timestamp 1636968456
transform 1 0 43148 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_152_469
timestamp 1
transform 1 0 44252 0 1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_152_475
timestamp 1
transform 1 0 44804 0 1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_152_477
timestamp 1636968456
transform 1 0 44988 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_489
timestamp 1636968456
transform 1 0 46092 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_501
timestamp 1636968456
transform 1 0 47196 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_513
timestamp 1636968456
transform 1 0 48300 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_152_525
timestamp 1
transform 1 0 49404 0 1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_152_531
timestamp 1
transform 1 0 49956 0 1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_152_533
timestamp 1636968456
transform 1 0 50140 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_545
timestamp 1636968456
transform 1 0 51244 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_557
timestamp 1636968456
transform 1 0 52348 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_569
timestamp 1636968456
transform 1 0 53452 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_152_581
timestamp 1
transform 1 0 54556 0 1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_152_587
timestamp 1
transform 1 0 55108 0 1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_152_589
timestamp 1636968456
transform 1 0 55292 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_601
timestamp 1636968456
transform 1 0 56396 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_613
timestamp 1636968456
transform 1 0 57500 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_625
timestamp 1636968456
transform 1 0 58604 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_152_637
timestamp 1
transform 1 0 59708 0 1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_152_643
timestamp 1
transform 1 0 60260 0 1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_152_645
timestamp 1636968456
transform 1 0 60444 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_657
timestamp 1636968456
transform 1 0 61548 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_669
timestamp 1636968456
transform 1 0 62652 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_681
timestamp 1636968456
transform 1 0 63756 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_152_693
timestamp 1
transform 1 0 64860 0 1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_152_699
timestamp 1
transform 1 0 65412 0 1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_152_701
timestamp 1636968456
transform 1 0 65596 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_713
timestamp 1636968456
transform 1 0 66700 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_725
timestamp 1636968456
transform 1 0 67804 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_737
timestamp 1636968456
transform 1 0 68908 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_152_749
timestamp 1
transform 1 0 70012 0 1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_152_755
timestamp 1
transform 1 0 70564 0 1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_152_757
timestamp 1636968456
transform 1 0 70748 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_769
timestamp 1636968456
transform 1 0 71852 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_781
timestamp 1636968456
transform 1 0 72956 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_793
timestamp 1636968456
transform 1 0 74060 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_152_805
timestamp 1
transform 1 0 75164 0 1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_152_811
timestamp 1
transform 1 0 75716 0 1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_152_813
timestamp 1636968456
transform 1 0 75900 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_825
timestamp 1636968456
transform 1 0 77004 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_837
timestamp 1636968456
transform 1 0 78108 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_849
timestamp 1636968456
transform 1 0 79212 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_152_861
timestamp 1
transform 1 0 80316 0 1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_152_867
timestamp 1
transform 1 0 80868 0 1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_152_869
timestamp 1636968456
transform 1 0 81052 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_881
timestamp 1636968456
transform 1 0 82156 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_893
timestamp 1636968456
transform 1 0 83260 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_905
timestamp 1636968456
transform 1 0 84364 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_152_917
timestamp 1
transform 1 0 85468 0 1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_152_923
timestamp 1
transform 1 0 86020 0 1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_152_925
timestamp 1636968456
transform 1 0 86204 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_937
timestamp 1636968456
transform 1 0 87308 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_949
timestamp 1636968456
transform 1 0 88412 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_961
timestamp 1636968456
transform 1 0 89516 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_152_973
timestamp 1
transform 1 0 90620 0 1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_152_979
timestamp 1
transform 1 0 91172 0 1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_152_981
timestamp 1636968456
transform 1 0 91356 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_993
timestamp 1636968456
transform 1 0 92460 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_1005
timestamp 1636968456
transform 1 0 93564 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_1017
timestamp 1636968456
transform 1 0 94668 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_152_1029
timestamp 1
transform 1 0 95772 0 1 84864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_152_1035
timestamp 1
transform 1 0 96324 0 1 84864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_152_1037
timestamp 1636968456
transform 1 0 96508 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_1049
timestamp 1636968456
transform 1 0 97612 0 1 84864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_1061
timestamp 1636968456
transform 1 0 98716 0 1 84864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_152_1073
timestamp 1
transform 1 0 99820 0 1 84864
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_153_3
timestamp 1636968456
transform 1 0 1380 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_15
timestamp 1636968456
transform 1 0 2484 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_27
timestamp 1636968456
transform 1 0 3588 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_39
timestamp 1636968456
transform 1 0 4692 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_153_51
timestamp 1
transform 1 0 5796 0 -1 85952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_153_55
timestamp 1
transform 1 0 6164 0 -1 85952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_153_57
timestamp 1636968456
transform 1 0 6348 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_69
timestamp 1636968456
transform 1 0 7452 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_81
timestamp 1636968456
transform 1 0 8556 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_93
timestamp 1636968456
transform 1 0 9660 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_153_105
timestamp 1
transform 1 0 10764 0 -1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_153_111
timestamp 1
transform 1 0 11316 0 -1 85952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_153_113
timestamp 1636968456
transform 1 0 11500 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_125
timestamp 1636968456
transform 1 0 12604 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_137
timestamp 1636968456
transform 1 0 13708 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_149
timestamp 1636968456
transform 1 0 14812 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_153_161
timestamp 1
transform 1 0 15916 0 -1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_153_167
timestamp 1
transform 1 0 16468 0 -1 85952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_153_169
timestamp 1636968456
transform 1 0 16652 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_181
timestamp 1636968456
transform 1 0 17756 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_193
timestamp 1636968456
transform 1 0 18860 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_205
timestamp 1636968456
transform 1 0 19964 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_153_217
timestamp 1
transform 1 0 21068 0 -1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_153_223
timestamp 1
transform 1 0 21620 0 -1 85952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_153_225
timestamp 1636968456
transform 1 0 21804 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_237
timestamp 1636968456
transform 1 0 22908 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_249
timestamp 1636968456
transform 1 0 24012 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_261
timestamp 1636968456
transform 1 0 25116 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_153_273
timestamp 1
transform 1 0 26220 0 -1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_153_279
timestamp 1
transform 1 0 26772 0 -1 85952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_153_281
timestamp 1636968456
transform 1 0 26956 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_293
timestamp 1636968456
transform 1 0 28060 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_305
timestamp 1636968456
transform 1 0 29164 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_317
timestamp 1636968456
transform 1 0 30268 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_153_329
timestamp 1
transform 1 0 31372 0 -1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_153_335
timestamp 1
transform 1 0 31924 0 -1 85952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_153_337
timestamp 1636968456
transform 1 0 32108 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_349
timestamp 1636968456
transform 1 0 33212 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_361
timestamp 1636968456
transform 1 0 34316 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_373
timestamp 1636968456
transform 1 0 35420 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_153_385
timestamp 1
transform 1 0 36524 0 -1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_153_391
timestamp 1
transform 1 0 37076 0 -1 85952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_153_393
timestamp 1636968456
transform 1 0 37260 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_405
timestamp 1636968456
transform 1 0 38364 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_417
timestamp 1636968456
transform 1 0 39468 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_429
timestamp 1636968456
transform 1 0 40572 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_153_441
timestamp 1
transform 1 0 41676 0 -1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_153_447
timestamp 1
transform 1 0 42228 0 -1 85952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_153_449
timestamp 1636968456
transform 1 0 42412 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_461
timestamp 1636968456
transform 1 0 43516 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_473
timestamp 1636968456
transform 1 0 44620 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_485
timestamp 1636968456
transform 1 0 45724 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_153_497
timestamp 1
transform 1 0 46828 0 -1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_153_503
timestamp 1
transform 1 0 47380 0 -1 85952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_153_505
timestamp 1636968456
transform 1 0 47564 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_517
timestamp 1636968456
transform 1 0 48668 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_529
timestamp 1636968456
transform 1 0 49772 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_541
timestamp 1636968456
transform 1 0 50876 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_153_553
timestamp 1
transform 1 0 51980 0 -1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_153_559
timestamp 1
transform 1 0 52532 0 -1 85952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_153_561
timestamp 1636968456
transform 1 0 52716 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_573
timestamp 1636968456
transform 1 0 53820 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_585
timestamp 1636968456
transform 1 0 54924 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_597
timestamp 1636968456
transform 1 0 56028 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_153_609
timestamp 1
transform 1 0 57132 0 -1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_153_615
timestamp 1
transform 1 0 57684 0 -1 85952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_153_617
timestamp 1636968456
transform 1 0 57868 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_629
timestamp 1636968456
transform 1 0 58972 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_641
timestamp 1636968456
transform 1 0 60076 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_653
timestamp 1636968456
transform 1 0 61180 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_153_665
timestamp 1
transform 1 0 62284 0 -1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_153_671
timestamp 1
transform 1 0 62836 0 -1 85952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_153_673
timestamp 1636968456
transform 1 0 63020 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_685
timestamp 1636968456
transform 1 0 64124 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_697
timestamp 1636968456
transform 1 0 65228 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_709
timestamp 1636968456
transform 1 0 66332 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_153_721
timestamp 1
transform 1 0 67436 0 -1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_153_727
timestamp 1
transform 1 0 67988 0 -1 85952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_153_729
timestamp 1636968456
transform 1 0 68172 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_741
timestamp 1636968456
transform 1 0 69276 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_753
timestamp 1636968456
transform 1 0 70380 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_765
timestamp 1636968456
transform 1 0 71484 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_153_777
timestamp 1
transform 1 0 72588 0 -1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_153_783
timestamp 1
transform 1 0 73140 0 -1 85952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_153_785
timestamp 1636968456
transform 1 0 73324 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_797
timestamp 1636968456
transform 1 0 74428 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_809
timestamp 1636968456
transform 1 0 75532 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_821
timestamp 1636968456
transform 1 0 76636 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_153_833
timestamp 1
transform 1 0 77740 0 -1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_153_839
timestamp 1
transform 1 0 78292 0 -1 85952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_153_841
timestamp 1636968456
transform 1 0 78476 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_853
timestamp 1636968456
transform 1 0 79580 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_865
timestamp 1636968456
transform 1 0 80684 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_877
timestamp 1636968456
transform 1 0 81788 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_153_889
timestamp 1
transform 1 0 82892 0 -1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_153_895
timestamp 1
transform 1 0 83444 0 -1 85952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_153_897
timestamp 1636968456
transform 1 0 83628 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_909
timestamp 1636968456
transform 1 0 84732 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_921
timestamp 1636968456
transform 1 0 85836 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_933
timestamp 1636968456
transform 1 0 86940 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_153_945
timestamp 1
transform 1 0 88044 0 -1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_153_951
timestamp 1
transform 1 0 88596 0 -1 85952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_153_953
timestamp 1636968456
transform 1 0 88780 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_965
timestamp 1636968456
transform 1 0 89884 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_977
timestamp 1636968456
transform 1 0 90988 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_989
timestamp 1636968456
transform 1 0 92092 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_153_1001
timestamp 1
transform 1 0 93196 0 -1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_153_1007
timestamp 1
transform 1 0 93748 0 -1 85952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_153_1009
timestamp 1636968456
transform 1 0 93932 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_1021
timestamp 1636968456
transform 1 0 95036 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_1033
timestamp 1636968456
transform 1 0 96140 0 -1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_1045
timestamp 1636968456
transform 1 0 97244 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_153_1057
timestamp 1
transform 1 0 98348 0 -1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_153_1063
timestamp 1
transform 1 0 98900 0 -1 85952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_153_1065
timestamp 1636968456
transform 1 0 99084 0 -1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_153_1077
timestamp 1
transform 1 0 100188 0 -1 85952
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_154_3
timestamp 1636968456
transform 1 0 1380 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_15
timestamp 1636968456
transform 1 0 2484 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_154_27
timestamp 1
transform 1 0 3588 0 1 85952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_154_29
timestamp 1636968456
transform 1 0 3772 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_41
timestamp 1636968456
transform 1 0 4876 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_53
timestamp 1636968456
transform 1 0 5980 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_65
timestamp 1636968456
transform 1 0 7084 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_154_77
timestamp 1
transform 1 0 8188 0 1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_154_83
timestamp 1
transform 1 0 8740 0 1 85952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_154_85
timestamp 1636968456
transform 1 0 8924 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_97
timestamp 1636968456
transform 1 0 10028 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_109
timestamp 1636968456
transform 1 0 11132 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_121
timestamp 1636968456
transform 1 0 12236 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_154_133
timestamp 1
transform 1 0 13340 0 1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_154_139
timestamp 1
transform 1 0 13892 0 1 85952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_154_141
timestamp 1636968456
transform 1 0 14076 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_153
timestamp 1636968456
transform 1 0 15180 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_165
timestamp 1636968456
transform 1 0 16284 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_177
timestamp 1636968456
transform 1 0 17388 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_154_189
timestamp 1
transform 1 0 18492 0 1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_154_195
timestamp 1
transform 1 0 19044 0 1 85952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_154_197
timestamp 1636968456
transform 1 0 19228 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_209
timestamp 1636968456
transform 1 0 20332 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_221
timestamp 1636968456
transform 1 0 21436 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_233
timestamp 1636968456
transform 1 0 22540 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_154_245
timestamp 1
transform 1 0 23644 0 1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_154_251
timestamp 1
transform 1 0 24196 0 1 85952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_154_253
timestamp 1636968456
transform 1 0 24380 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_265
timestamp 1636968456
transform 1 0 25484 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_277
timestamp 1636968456
transform 1 0 26588 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_289
timestamp 1636968456
transform 1 0 27692 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_154_301
timestamp 1
transform 1 0 28796 0 1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_154_307
timestamp 1
transform 1 0 29348 0 1 85952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_154_309
timestamp 1636968456
transform 1 0 29532 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_321
timestamp 1636968456
transform 1 0 30636 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_333
timestamp 1636968456
transform 1 0 31740 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_345
timestamp 1636968456
transform 1 0 32844 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_154_357
timestamp 1
transform 1 0 33948 0 1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_154_363
timestamp 1
transform 1 0 34500 0 1 85952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_154_365
timestamp 1636968456
transform 1 0 34684 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_377
timestamp 1636968456
transform 1 0 35788 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_389
timestamp 1636968456
transform 1 0 36892 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_401
timestamp 1636968456
transform 1 0 37996 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_154_413
timestamp 1
transform 1 0 39100 0 1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_154_419
timestamp 1
transform 1 0 39652 0 1 85952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_154_421
timestamp 1636968456
transform 1 0 39836 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_433
timestamp 1636968456
transform 1 0 40940 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_445
timestamp 1636968456
transform 1 0 42044 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_457
timestamp 1636968456
transform 1 0 43148 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_154_469
timestamp 1
transform 1 0 44252 0 1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_154_475
timestamp 1
transform 1 0 44804 0 1 85952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_154_477
timestamp 1636968456
transform 1 0 44988 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_489
timestamp 1636968456
transform 1 0 46092 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_501
timestamp 1636968456
transform 1 0 47196 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_513
timestamp 1636968456
transform 1 0 48300 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_154_525
timestamp 1
transform 1 0 49404 0 1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_154_531
timestamp 1
transform 1 0 49956 0 1 85952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_154_533
timestamp 1636968456
transform 1 0 50140 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_545
timestamp 1636968456
transform 1 0 51244 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_557
timestamp 1636968456
transform 1 0 52348 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_569
timestamp 1636968456
transform 1 0 53452 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_154_581
timestamp 1
transform 1 0 54556 0 1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_154_587
timestamp 1
transform 1 0 55108 0 1 85952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_154_589
timestamp 1636968456
transform 1 0 55292 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_601
timestamp 1636968456
transform 1 0 56396 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_613
timestamp 1636968456
transform 1 0 57500 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_625
timestamp 1636968456
transform 1 0 58604 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_154_637
timestamp 1
transform 1 0 59708 0 1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_154_643
timestamp 1
transform 1 0 60260 0 1 85952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_154_645
timestamp 1636968456
transform 1 0 60444 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_657
timestamp 1636968456
transform 1 0 61548 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_669
timestamp 1636968456
transform 1 0 62652 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_681
timestamp 1636968456
transform 1 0 63756 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_154_693
timestamp 1
transform 1 0 64860 0 1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_154_699
timestamp 1
transform 1 0 65412 0 1 85952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_154_701
timestamp 1636968456
transform 1 0 65596 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_713
timestamp 1636968456
transform 1 0 66700 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_725
timestamp 1636968456
transform 1 0 67804 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_737
timestamp 1636968456
transform 1 0 68908 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_154_749
timestamp 1
transform 1 0 70012 0 1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_154_755
timestamp 1
transform 1 0 70564 0 1 85952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_154_757
timestamp 1636968456
transform 1 0 70748 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_769
timestamp 1636968456
transform 1 0 71852 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_781
timestamp 1636968456
transform 1 0 72956 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_793
timestamp 1636968456
transform 1 0 74060 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_154_805
timestamp 1
transform 1 0 75164 0 1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_154_811
timestamp 1
transform 1 0 75716 0 1 85952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_154_813
timestamp 1636968456
transform 1 0 75900 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_825
timestamp 1636968456
transform 1 0 77004 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_837
timestamp 1636968456
transform 1 0 78108 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_849
timestamp 1636968456
transform 1 0 79212 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_154_861
timestamp 1
transform 1 0 80316 0 1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_154_867
timestamp 1
transform 1 0 80868 0 1 85952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_154_869
timestamp 1636968456
transform 1 0 81052 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_881
timestamp 1636968456
transform 1 0 82156 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_893
timestamp 1636968456
transform 1 0 83260 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_905
timestamp 1636968456
transform 1 0 84364 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_154_917
timestamp 1
transform 1 0 85468 0 1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_154_923
timestamp 1
transform 1 0 86020 0 1 85952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_154_925
timestamp 1636968456
transform 1 0 86204 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_937
timestamp 1636968456
transform 1 0 87308 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_949
timestamp 1636968456
transform 1 0 88412 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_961
timestamp 1636968456
transform 1 0 89516 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_154_973
timestamp 1
transform 1 0 90620 0 1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_154_979
timestamp 1
transform 1 0 91172 0 1 85952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_154_981
timestamp 1636968456
transform 1 0 91356 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_993
timestamp 1636968456
transform 1 0 92460 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_1005
timestamp 1636968456
transform 1 0 93564 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_1017
timestamp 1636968456
transform 1 0 94668 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_154_1029
timestamp 1
transform 1 0 95772 0 1 85952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_154_1035
timestamp 1
transform 1 0 96324 0 1 85952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_154_1037
timestamp 1636968456
transform 1 0 96508 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_1049
timestamp 1636968456
transform 1 0 97612 0 1 85952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_1061
timestamp 1636968456
transform 1 0 98716 0 1 85952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_154_1073
timestamp 1
transform 1 0 99820 0 1 85952
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_155_3
timestamp 1636968456
transform 1 0 1380 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_15
timestamp 1636968456
transform 1 0 2484 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_27
timestamp 1636968456
transform 1 0 3588 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_39
timestamp 1636968456
transform 1 0 4692 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_155_51
timestamp 1
transform 1 0 5796 0 -1 87040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_155_55
timestamp 1
transform 1 0 6164 0 -1 87040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_155_57
timestamp 1636968456
transform 1 0 6348 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_69
timestamp 1636968456
transform 1 0 7452 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_81
timestamp 1636968456
transform 1 0 8556 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_93
timestamp 1636968456
transform 1 0 9660 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_155_105
timestamp 1
transform 1 0 10764 0 -1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_155_111
timestamp 1
transform 1 0 11316 0 -1 87040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_155_113
timestamp 1636968456
transform 1 0 11500 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_125
timestamp 1636968456
transform 1 0 12604 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_137
timestamp 1636968456
transform 1 0 13708 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_149
timestamp 1636968456
transform 1 0 14812 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_155_161
timestamp 1
transform 1 0 15916 0 -1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_155_167
timestamp 1
transform 1 0 16468 0 -1 87040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_155_169
timestamp 1636968456
transform 1 0 16652 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_181
timestamp 1636968456
transform 1 0 17756 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_193
timestamp 1636968456
transform 1 0 18860 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_205
timestamp 1636968456
transform 1 0 19964 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_155_217
timestamp 1
transform 1 0 21068 0 -1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_155_223
timestamp 1
transform 1 0 21620 0 -1 87040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_155_225
timestamp 1636968456
transform 1 0 21804 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_237
timestamp 1636968456
transform 1 0 22908 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_249
timestamp 1636968456
transform 1 0 24012 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_261
timestamp 1636968456
transform 1 0 25116 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_155_273
timestamp 1
transform 1 0 26220 0 -1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_155_279
timestamp 1
transform 1 0 26772 0 -1 87040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_155_281
timestamp 1636968456
transform 1 0 26956 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_293
timestamp 1636968456
transform 1 0 28060 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_305
timestamp 1636968456
transform 1 0 29164 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_317
timestamp 1636968456
transform 1 0 30268 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_155_329
timestamp 1
transform 1 0 31372 0 -1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_155_335
timestamp 1
transform 1 0 31924 0 -1 87040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_155_337
timestamp 1636968456
transform 1 0 32108 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_349
timestamp 1636968456
transform 1 0 33212 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_361
timestamp 1636968456
transform 1 0 34316 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_373
timestamp 1636968456
transform 1 0 35420 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_155_385
timestamp 1
transform 1 0 36524 0 -1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_155_391
timestamp 1
transform 1 0 37076 0 -1 87040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_155_393
timestamp 1636968456
transform 1 0 37260 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_405
timestamp 1636968456
transform 1 0 38364 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_417
timestamp 1636968456
transform 1 0 39468 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_429
timestamp 1636968456
transform 1 0 40572 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_155_441
timestamp 1
transform 1 0 41676 0 -1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_155_447
timestamp 1
transform 1 0 42228 0 -1 87040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_155_449
timestamp 1636968456
transform 1 0 42412 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_461
timestamp 1636968456
transform 1 0 43516 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_473
timestamp 1636968456
transform 1 0 44620 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_485
timestamp 1636968456
transform 1 0 45724 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_155_497
timestamp 1
transform 1 0 46828 0 -1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_155_503
timestamp 1
transform 1 0 47380 0 -1 87040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_155_505
timestamp 1636968456
transform 1 0 47564 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_517
timestamp 1636968456
transform 1 0 48668 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_529
timestamp 1636968456
transform 1 0 49772 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_541
timestamp 1636968456
transform 1 0 50876 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_155_553
timestamp 1
transform 1 0 51980 0 -1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_155_559
timestamp 1
transform 1 0 52532 0 -1 87040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_155_561
timestamp 1636968456
transform 1 0 52716 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_573
timestamp 1636968456
transform 1 0 53820 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_585
timestamp 1636968456
transform 1 0 54924 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_597
timestamp 1636968456
transform 1 0 56028 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_155_609
timestamp 1
transform 1 0 57132 0 -1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_155_615
timestamp 1
transform 1 0 57684 0 -1 87040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_155_617
timestamp 1636968456
transform 1 0 57868 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_629
timestamp 1636968456
transform 1 0 58972 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_641
timestamp 1636968456
transform 1 0 60076 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_653
timestamp 1636968456
transform 1 0 61180 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_155_665
timestamp 1
transform 1 0 62284 0 -1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_155_671
timestamp 1
transform 1 0 62836 0 -1 87040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_155_673
timestamp 1636968456
transform 1 0 63020 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_685
timestamp 1636968456
transform 1 0 64124 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_697
timestamp 1636968456
transform 1 0 65228 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_709
timestamp 1636968456
transform 1 0 66332 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_155_721
timestamp 1
transform 1 0 67436 0 -1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_155_727
timestamp 1
transform 1 0 67988 0 -1 87040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_155_729
timestamp 1636968456
transform 1 0 68172 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_741
timestamp 1636968456
transform 1 0 69276 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_753
timestamp 1636968456
transform 1 0 70380 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_765
timestamp 1636968456
transform 1 0 71484 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_155_777
timestamp 1
transform 1 0 72588 0 -1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_155_783
timestamp 1
transform 1 0 73140 0 -1 87040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_155_785
timestamp 1636968456
transform 1 0 73324 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_797
timestamp 1636968456
transform 1 0 74428 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_809
timestamp 1636968456
transform 1 0 75532 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_821
timestamp 1636968456
transform 1 0 76636 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_155_833
timestamp 1
transform 1 0 77740 0 -1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_155_839
timestamp 1
transform 1 0 78292 0 -1 87040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_155_841
timestamp 1636968456
transform 1 0 78476 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_853
timestamp 1636968456
transform 1 0 79580 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_865
timestamp 1636968456
transform 1 0 80684 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_877
timestamp 1636968456
transform 1 0 81788 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_155_889
timestamp 1
transform 1 0 82892 0 -1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_155_895
timestamp 1
transform 1 0 83444 0 -1 87040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_155_897
timestamp 1636968456
transform 1 0 83628 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_909
timestamp 1636968456
transform 1 0 84732 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_921
timestamp 1636968456
transform 1 0 85836 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_933
timestamp 1636968456
transform 1 0 86940 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_155_945
timestamp 1
transform 1 0 88044 0 -1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_155_951
timestamp 1
transform 1 0 88596 0 -1 87040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_155_953
timestamp 1636968456
transform 1 0 88780 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_965
timestamp 1636968456
transform 1 0 89884 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_977
timestamp 1636968456
transform 1 0 90988 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_989
timestamp 1636968456
transform 1 0 92092 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_155_1001
timestamp 1
transform 1 0 93196 0 -1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_155_1007
timestamp 1
transform 1 0 93748 0 -1 87040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_155_1009
timestamp 1636968456
transform 1 0 93932 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_1021
timestamp 1636968456
transform 1 0 95036 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_1033
timestamp 1636968456
transform 1 0 96140 0 -1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_155_1045
timestamp 1636968456
transform 1 0 97244 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_155_1057
timestamp 1
transform 1 0 98348 0 -1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_155_1063
timestamp 1
transform 1 0 98900 0 -1 87040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_155_1065
timestamp 1636968456
transform 1 0 99084 0 -1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_155_1077
timestamp 1
transform 1 0 100188 0 -1 87040
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_156_3
timestamp 1636968456
transform 1 0 1380 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_15
timestamp 1636968456
transform 1 0 2484 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_156_27
timestamp 1
transform 1 0 3588 0 1 87040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_156_29
timestamp 1636968456
transform 1 0 3772 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_41
timestamp 1636968456
transform 1 0 4876 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_53
timestamp 1636968456
transform 1 0 5980 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_65
timestamp 1636968456
transform 1 0 7084 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_156_77
timestamp 1
transform 1 0 8188 0 1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_156_83
timestamp 1
transform 1 0 8740 0 1 87040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_156_85
timestamp 1636968456
transform 1 0 8924 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_97
timestamp 1636968456
transform 1 0 10028 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_109
timestamp 1636968456
transform 1 0 11132 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_121
timestamp 1636968456
transform 1 0 12236 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_156_133
timestamp 1
transform 1 0 13340 0 1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_156_139
timestamp 1
transform 1 0 13892 0 1 87040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_156_141
timestamp 1636968456
transform 1 0 14076 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_153
timestamp 1636968456
transform 1 0 15180 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_165
timestamp 1636968456
transform 1 0 16284 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_177
timestamp 1636968456
transform 1 0 17388 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_156_189
timestamp 1
transform 1 0 18492 0 1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_156_195
timestamp 1
transform 1 0 19044 0 1 87040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_156_197
timestamp 1636968456
transform 1 0 19228 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_209
timestamp 1636968456
transform 1 0 20332 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_221
timestamp 1636968456
transform 1 0 21436 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_233
timestamp 1636968456
transform 1 0 22540 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_156_245
timestamp 1
transform 1 0 23644 0 1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_156_251
timestamp 1
transform 1 0 24196 0 1 87040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_156_253
timestamp 1636968456
transform 1 0 24380 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_265
timestamp 1636968456
transform 1 0 25484 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_277
timestamp 1636968456
transform 1 0 26588 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_289
timestamp 1636968456
transform 1 0 27692 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_156_301
timestamp 1
transform 1 0 28796 0 1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_156_307
timestamp 1
transform 1 0 29348 0 1 87040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_156_309
timestamp 1636968456
transform 1 0 29532 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_321
timestamp 1636968456
transform 1 0 30636 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_333
timestamp 1636968456
transform 1 0 31740 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_345
timestamp 1636968456
transform 1 0 32844 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_156_357
timestamp 1
transform 1 0 33948 0 1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_156_363
timestamp 1
transform 1 0 34500 0 1 87040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_156_365
timestamp 1636968456
transform 1 0 34684 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_377
timestamp 1636968456
transform 1 0 35788 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_389
timestamp 1636968456
transform 1 0 36892 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_401
timestamp 1636968456
transform 1 0 37996 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_156_413
timestamp 1
transform 1 0 39100 0 1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_156_419
timestamp 1
transform 1 0 39652 0 1 87040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_156_421
timestamp 1636968456
transform 1 0 39836 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_433
timestamp 1636968456
transform 1 0 40940 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_445
timestamp 1636968456
transform 1 0 42044 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_457
timestamp 1636968456
transform 1 0 43148 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_156_469
timestamp 1
transform 1 0 44252 0 1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_156_475
timestamp 1
transform 1 0 44804 0 1 87040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_156_477
timestamp 1636968456
transform 1 0 44988 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_489
timestamp 1636968456
transform 1 0 46092 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_501
timestamp 1636968456
transform 1 0 47196 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_513
timestamp 1636968456
transform 1 0 48300 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_156_525
timestamp 1
transform 1 0 49404 0 1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_156_531
timestamp 1
transform 1 0 49956 0 1 87040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_156_533
timestamp 1636968456
transform 1 0 50140 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_545
timestamp 1636968456
transform 1 0 51244 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_557
timestamp 1636968456
transform 1 0 52348 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_569
timestamp 1636968456
transform 1 0 53452 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_156_581
timestamp 1
transform 1 0 54556 0 1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_156_587
timestamp 1
transform 1 0 55108 0 1 87040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_156_589
timestamp 1636968456
transform 1 0 55292 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_601
timestamp 1636968456
transform 1 0 56396 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_613
timestamp 1636968456
transform 1 0 57500 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_625
timestamp 1636968456
transform 1 0 58604 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_156_637
timestamp 1
transform 1 0 59708 0 1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_156_643
timestamp 1
transform 1 0 60260 0 1 87040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_156_645
timestamp 1636968456
transform 1 0 60444 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_657
timestamp 1636968456
transform 1 0 61548 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_669
timestamp 1636968456
transform 1 0 62652 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_681
timestamp 1636968456
transform 1 0 63756 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_156_693
timestamp 1
transform 1 0 64860 0 1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_156_699
timestamp 1
transform 1 0 65412 0 1 87040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_156_701
timestamp 1636968456
transform 1 0 65596 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_713
timestamp 1636968456
transform 1 0 66700 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_725
timestamp 1636968456
transform 1 0 67804 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_737
timestamp 1636968456
transform 1 0 68908 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_156_749
timestamp 1
transform 1 0 70012 0 1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_156_755
timestamp 1
transform 1 0 70564 0 1 87040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_156_757
timestamp 1636968456
transform 1 0 70748 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_769
timestamp 1636968456
transform 1 0 71852 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_781
timestamp 1636968456
transform 1 0 72956 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_793
timestamp 1636968456
transform 1 0 74060 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_156_805
timestamp 1
transform 1 0 75164 0 1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_156_811
timestamp 1
transform 1 0 75716 0 1 87040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_156_813
timestamp 1636968456
transform 1 0 75900 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_825
timestamp 1636968456
transform 1 0 77004 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_837
timestamp 1636968456
transform 1 0 78108 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_849
timestamp 1636968456
transform 1 0 79212 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_156_861
timestamp 1
transform 1 0 80316 0 1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_156_867
timestamp 1
transform 1 0 80868 0 1 87040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_156_869
timestamp 1636968456
transform 1 0 81052 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_881
timestamp 1636968456
transform 1 0 82156 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_893
timestamp 1636968456
transform 1 0 83260 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_905
timestamp 1636968456
transform 1 0 84364 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_156_917
timestamp 1
transform 1 0 85468 0 1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_156_923
timestamp 1
transform 1 0 86020 0 1 87040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_156_925
timestamp 1636968456
transform 1 0 86204 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_937
timestamp 1636968456
transform 1 0 87308 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_949
timestamp 1636968456
transform 1 0 88412 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_961
timestamp 1636968456
transform 1 0 89516 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_156_973
timestamp 1
transform 1 0 90620 0 1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_156_979
timestamp 1
transform 1 0 91172 0 1 87040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_156_981
timestamp 1636968456
transform 1 0 91356 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_993
timestamp 1636968456
transform 1 0 92460 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_1005
timestamp 1636968456
transform 1 0 93564 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_1017
timestamp 1636968456
transform 1 0 94668 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_156_1029
timestamp 1
transform 1 0 95772 0 1 87040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_156_1035
timestamp 1
transform 1 0 96324 0 1 87040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_156_1037
timestamp 1636968456
transform 1 0 96508 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_1049
timestamp 1636968456
transform 1 0 97612 0 1 87040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_156_1061
timestamp 1636968456
transform 1 0 98716 0 1 87040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_156_1073
timestamp 1
transform 1 0 99820 0 1 87040
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_157_3
timestamp 1636968456
transform 1 0 1380 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_15
timestamp 1636968456
transform 1 0 2484 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_27
timestamp 1636968456
transform 1 0 3588 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_39
timestamp 1636968456
transform 1 0 4692 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_157_51
timestamp 1
transform 1 0 5796 0 -1 88128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_157_55
timestamp 1
transform 1 0 6164 0 -1 88128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_157_57
timestamp 1636968456
transform 1 0 6348 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_69
timestamp 1636968456
transform 1 0 7452 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_81
timestamp 1636968456
transform 1 0 8556 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_93
timestamp 1636968456
transform 1 0 9660 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_157_105
timestamp 1
transform 1 0 10764 0 -1 88128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_157_111
timestamp 1
transform 1 0 11316 0 -1 88128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_157_113
timestamp 1636968456
transform 1 0 11500 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_125
timestamp 1636968456
transform 1 0 12604 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_137
timestamp 1636968456
transform 1 0 13708 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_149
timestamp 1636968456
transform 1 0 14812 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_157_161
timestamp 1
transform 1 0 15916 0 -1 88128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_157_167
timestamp 1
transform 1 0 16468 0 -1 88128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_157_169
timestamp 1636968456
transform 1 0 16652 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_181
timestamp 1636968456
transform 1 0 17756 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_193
timestamp 1636968456
transform 1 0 18860 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_205
timestamp 1636968456
transform 1 0 19964 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_157_217
timestamp 1
transform 1 0 21068 0 -1 88128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_157_223
timestamp 1
transform 1 0 21620 0 -1 88128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_157_225
timestamp 1636968456
transform 1 0 21804 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_237
timestamp 1636968456
transform 1 0 22908 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_249
timestamp 1636968456
transform 1 0 24012 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_261
timestamp 1636968456
transform 1 0 25116 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_157_273
timestamp 1
transform 1 0 26220 0 -1 88128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_157_279
timestamp 1
transform 1 0 26772 0 -1 88128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_157_281
timestamp 1636968456
transform 1 0 26956 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_293
timestamp 1636968456
transform 1 0 28060 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_305
timestamp 1636968456
transform 1 0 29164 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_317
timestamp 1636968456
transform 1 0 30268 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_157_329
timestamp 1
transform 1 0 31372 0 -1 88128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_157_335
timestamp 1
transform 1 0 31924 0 -1 88128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_157_337
timestamp 1636968456
transform 1 0 32108 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_349
timestamp 1636968456
transform 1 0 33212 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_361
timestamp 1636968456
transform 1 0 34316 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_373
timestamp 1636968456
transform 1 0 35420 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_157_385
timestamp 1
transform 1 0 36524 0 -1 88128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_157_391
timestamp 1
transform 1 0 37076 0 -1 88128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_157_393
timestamp 1636968456
transform 1 0 37260 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_405
timestamp 1636968456
transform 1 0 38364 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_417
timestamp 1636968456
transform 1 0 39468 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_429
timestamp 1636968456
transform 1 0 40572 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_157_441
timestamp 1
transform 1 0 41676 0 -1 88128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_157_447
timestamp 1
transform 1 0 42228 0 -1 88128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_157_449
timestamp 1636968456
transform 1 0 42412 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_461
timestamp 1636968456
transform 1 0 43516 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_473
timestamp 1636968456
transform 1 0 44620 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_485
timestamp 1636968456
transform 1 0 45724 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_157_497
timestamp 1
transform 1 0 46828 0 -1 88128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_157_503
timestamp 1
transform 1 0 47380 0 -1 88128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_157_505
timestamp 1636968456
transform 1 0 47564 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_517
timestamp 1636968456
transform 1 0 48668 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_529
timestamp 1636968456
transform 1 0 49772 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_541
timestamp 1636968456
transform 1 0 50876 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_157_553
timestamp 1
transform 1 0 51980 0 -1 88128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_157_559
timestamp 1
transform 1 0 52532 0 -1 88128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_157_561
timestamp 1636968456
transform 1 0 52716 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_573
timestamp 1636968456
transform 1 0 53820 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_585
timestamp 1636968456
transform 1 0 54924 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_597
timestamp 1636968456
transform 1 0 56028 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_157_609
timestamp 1
transform 1 0 57132 0 -1 88128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_157_615
timestamp 1
transform 1 0 57684 0 -1 88128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_157_617
timestamp 1636968456
transform 1 0 57868 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_629
timestamp 1636968456
transform 1 0 58972 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_641
timestamp 1636968456
transform 1 0 60076 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_653
timestamp 1636968456
transform 1 0 61180 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_157_665
timestamp 1
transform 1 0 62284 0 -1 88128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_157_671
timestamp 1
transform 1 0 62836 0 -1 88128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_157_673
timestamp 1636968456
transform 1 0 63020 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_685
timestamp 1636968456
transform 1 0 64124 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_697
timestamp 1636968456
transform 1 0 65228 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_709
timestamp 1636968456
transform 1 0 66332 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_157_721
timestamp 1
transform 1 0 67436 0 -1 88128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_157_727
timestamp 1
transform 1 0 67988 0 -1 88128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_157_729
timestamp 1636968456
transform 1 0 68172 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_741
timestamp 1636968456
transform 1 0 69276 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_753
timestamp 1636968456
transform 1 0 70380 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_765
timestamp 1636968456
transform 1 0 71484 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_157_777
timestamp 1
transform 1 0 72588 0 -1 88128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_157_783
timestamp 1
transform 1 0 73140 0 -1 88128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_157_785
timestamp 1636968456
transform 1 0 73324 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_797
timestamp 1636968456
transform 1 0 74428 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_809
timestamp 1636968456
transform 1 0 75532 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_821
timestamp 1636968456
transform 1 0 76636 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_157_833
timestamp 1
transform 1 0 77740 0 -1 88128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_157_839
timestamp 1
transform 1 0 78292 0 -1 88128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_157_841
timestamp 1636968456
transform 1 0 78476 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_853
timestamp 1636968456
transform 1 0 79580 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_865
timestamp 1636968456
transform 1 0 80684 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_877
timestamp 1636968456
transform 1 0 81788 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_157_889
timestamp 1
transform 1 0 82892 0 -1 88128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_157_895
timestamp 1
transform 1 0 83444 0 -1 88128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_157_897
timestamp 1636968456
transform 1 0 83628 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_909
timestamp 1636968456
transform 1 0 84732 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_921
timestamp 1636968456
transform 1 0 85836 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_933
timestamp 1636968456
transform 1 0 86940 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_157_945
timestamp 1
transform 1 0 88044 0 -1 88128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_157_951
timestamp 1
transform 1 0 88596 0 -1 88128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_157_953
timestamp 1636968456
transform 1 0 88780 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_965
timestamp 1636968456
transform 1 0 89884 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_977
timestamp 1636968456
transform 1 0 90988 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_989
timestamp 1636968456
transform 1 0 92092 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_157_1001
timestamp 1
transform 1 0 93196 0 -1 88128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_157_1007
timestamp 1
transform 1 0 93748 0 -1 88128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_157_1009
timestamp 1636968456
transform 1 0 93932 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_1021
timestamp 1636968456
transform 1 0 95036 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_1033
timestamp 1636968456
transform 1 0 96140 0 -1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_157_1045
timestamp 1636968456
transform 1 0 97244 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_157_1057
timestamp 1
transform 1 0 98348 0 -1 88128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_157_1063
timestamp 1
transform 1 0 98900 0 -1 88128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_157_1065
timestamp 1636968456
transform 1 0 99084 0 -1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_157_1077
timestamp 1
transform 1 0 100188 0 -1 88128
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_158_3
timestamp 1636968456
transform 1 0 1380 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_15
timestamp 1636968456
transform 1 0 2484 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_158_27
timestamp 1
transform 1 0 3588 0 1 88128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_158_29
timestamp 1636968456
transform 1 0 3772 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_41
timestamp 1636968456
transform 1 0 4876 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_53
timestamp 1636968456
transform 1 0 5980 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_65
timestamp 1636968456
transform 1 0 7084 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_158_77
timestamp 1
transform 1 0 8188 0 1 88128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_158_83
timestamp 1
transform 1 0 8740 0 1 88128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_158_85
timestamp 1636968456
transform 1 0 8924 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_97
timestamp 1636968456
transform 1 0 10028 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_109
timestamp 1636968456
transform 1 0 11132 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_121
timestamp 1636968456
transform 1 0 12236 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_158_133
timestamp 1
transform 1 0 13340 0 1 88128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_158_139
timestamp 1
transform 1 0 13892 0 1 88128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_158_141
timestamp 1636968456
transform 1 0 14076 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_153
timestamp 1636968456
transform 1 0 15180 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_165
timestamp 1636968456
transform 1 0 16284 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_177
timestamp 1636968456
transform 1 0 17388 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_158_189
timestamp 1
transform 1 0 18492 0 1 88128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_158_195
timestamp 1
transform 1 0 19044 0 1 88128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_158_197
timestamp 1636968456
transform 1 0 19228 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_209
timestamp 1636968456
transform 1 0 20332 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_221
timestamp 1636968456
transform 1 0 21436 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_233
timestamp 1636968456
transform 1 0 22540 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_158_245
timestamp 1
transform 1 0 23644 0 1 88128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_158_251
timestamp 1
transform 1 0 24196 0 1 88128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_158_253
timestamp 1636968456
transform 1 0 24380 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_265
timestamp 1636968456
transform 1 0 25484 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_277
timestamp 1636968456
transform 1 0 26588 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_289
timestamp 1636968456
transform 1 0 27692 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_158_301
timestamp 1
transform 1 0 28796 0 1 88128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_158_307
timestamp 1
transform 1 0 29348 0 1 88128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_158_309
timestamp 1636968456
transform 1 0 29532 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_321
timestamp 1636968456
transform 1 0 30636 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_333
timestamp 1636968456
transform 1 0 31740 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_345
timestamp 1636968456
transform 1 0 32844 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_158_357
timestamp 1
transform 1 0 33948 0 1 88128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_158_363
timestamp 1
transform 1 0 34500 0 1 88128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_158_365
timestamp 1636968456
transform 1 0 34684 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_377
timestamp 1636968456
transform 1 0 35788 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_389
timestamp 1636968456
transform 1 0 36892 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_401
timestamp 1636968456
transform 1 0 37996 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_158_413
timestamp 1
transform 1 0 39100 0 1 88128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_158_419
timestamp 1
transform 1 0 39652 0 1 88128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_158_421
timestamp 1636968456
transform 1 0 39836 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_433
timestamp 1636968456
transform 1 0 40940 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_445
timestamp 1636968456
transform 1 0 42044 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_457
timestamp 1636968456
transform 1 0 43148 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_158_469
timestamp 1
transform 1 0 44252 0 1 88128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_158_475
timestamp 1
transform 1 0 44804 0 1 88128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_158_477
timestamp 1636968456
transform 1 0 44988 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_489
timestamp 1636968456
transform 1 0 46092 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_501
timestamp 1636968456
transform 1 0 47196 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_513
timestamp 1636968456
transform 1 0 48300 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_158_525
timestamp 1
transform 1 0 49404 0 1 88128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_158_531
timestamp 1
transform 1 0 49956 0 1 88128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_158_533
timestamp 1636968456
transform 1 0 50140 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_545
timestamp 1636968456
transform 1 0 51244 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_557
timestamp 1636968456
transform 1 0 52348 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_569
timestamp 1636968456
transform 1 0 53452 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_158_581
timestamp 1
transform 1 0 54556 0 1 88128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_158_587
timestamp 1
transform 1 0 55108 0 1 88128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_158_589
timestamp 1636968456
transform 1 0 55292 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_601
timestamp 1636968456
transform 1 0 56396 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_613
timestamp 1636968456
transform 1 0 57500 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_625
timestamp 1636968456
transform 1 0 58604 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_158_637
timestamp 1
transform 1 0 59708 0 1 88128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_158_643
timestamp 1
transform 1 0 60260 0 1 88128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_158_645
timestamp 1636968456
transform 1 0 60444 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_657
timestamp 1636968456
transform 1 0 61548 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_669
timestamp 1636968456
transform 1 0 62652 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_681
timestamp 1636968456
transform 1 0 63756 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_158_693
timestamp 1
transform 1 0 64860 0 1 88128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_158_699
timestamp 1
transform 1 0 65412 0 1 88128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_158_701
timestamp 1636968456
transform 1 0 65596 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_713
timestamp 1636968456
transform 1 0 66700 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_725
timestamp 1636968456
transform 1 0 67804 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_737
timestamp 1636968456
transform 1 0 68908 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_158_749
timestamp 1
transform 1 0 70012 0 1 88128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_158_755
timestamp 1
transform 1 0 70564 0 1 88128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_158_757
timestamp 1636968456
transform 1 0 70748 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_769
timestamp 1636968456
transform 1 0 71852 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_781
timestamp 1636968456
transform 1 0 72956 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_793
timestamp 1636968456
transform 1 0 74060 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_158_805
timestamp 1
transform 1 0 75164 0 1 88128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_158_811
timestamp 1
transform 1 0 75716 0 1 88128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_158_813
timestamp 1636968456
transform 1 0 75900 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_825
timestamp 1636968456
transform 1 0 77004 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_837
timestamp 1636968456
transform 1 0 78108 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_849
timestamp 1636968456
transform 1 0 79212 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_158_861
timestamp 1
transform 1 0 80316 0 1 88128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_158_867
timestamp 1
transform 1 0 80868 0 1 88128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_158_869
timestamp 1636968456
transform 1 0 81052 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_881
timestamp 1636968456
transform 1 0 82156 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_893
timestamp 1636968456
transform 1 0 83260 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_905
timestamp 1636968456
transform 1 0 84364 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_158_917
timestamp 1
transform 1 0 85468 0 1 88128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_158_923
timestamp 1
transform 1 0 86020 0 1 88128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_158_925
timestamp 1636968456
transform 1 0 86204 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_937
timestamp 1636968456
transform 1 0 87308 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_949
timestamp 1636968456
transform 1 0 88412 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_961
timestamp 1636968456
transform 1 0 89516 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_158_973
timestamp 1
transform 1 0 90620 0 1 88128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_158_979
timestamp 1
transform 1 0 91172 0 1 88128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_158_981
timestamp 1636968456
transform 1 0 91356 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_993
timestamp 1636968456
transform 1 0 92460 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_1005
timestamp 1636968456
transform 1 0 93564 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_1017
timestamp 1636968456
transform 1 0 94668 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_158_1029
timestamp 1
transform 1 0 95772 0 1 88128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_158_1035
timestamp 1
transform 1 0 96324 0 1 88128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_158_1037
timestamp 1636968456
transform 1 0 96508 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_1049
timestamp 1636968456
transform 1 0 97612 0 1 88128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_158_1061
timestamp 1636968456
transform 1 0 98716 0 1 88128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_158_1073
timestamp 1
transform 1 0 99820 0 1 88128
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_159_3
timestamp 1636968456
transform 1 0 1380 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_15
timestamp 1636968456
transform 1 0 2484 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_27
timestamp 1636968456
transform 1 0 3588 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_39
timestamp 1636968456
transform 1 0 4692 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_159_51
timestamp 1
transform 1 0 5796 0 -1 89216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_159_55
timestamp 1
transform 1 0 6164 0 -1 89216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_159_57
timestamp 1636968456
transform 1 0 6348 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_69
timestamp 1636968456
transform 1 0 7452 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_81
timestamp 1636968456
transform 1 0 8556 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_93
timestamp 1636968456
transform 1 0 9660 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_159_105
timestamp 1
transform 1 0 10764 0 -1 89216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_159_111
timestamp 1
transform 1 0 11316 0 -1 89216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_159_113
timestamp 1636968456
transform 1 0 11500 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_125
timestamp 1636968456
transform 1 0 12604 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_137
timestamp 1636968456
transform 1 0 13708 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_149
timestamp 1636968456
transform 1 0 14812 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_159_161
timestamp 1
transform 1 0 15916 0 -1 89216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_159_167
timestamp 1
transform 1 0 16468 0 -1 89216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_159_169
timestamp 1636968456
transform 1 0 16652 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_181
timestamp 1636968456
transform 1 0 17756 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_193
timestamp 1636968456
transform 1 0 18860 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_205
timestamp 1636968456
transform 1 0 19964 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_159_217
timestamp 1
transform 1 0 21068 0 -1 89216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_159_223
timestamp 1
transform 1 0 21620 0 -1 89216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_159_225
timestamp 1636968456
transform 1 0 21804 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_237
timestamp 1636968456
transform 1 0 22908 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_249
timestamp 1636968456
transform 1 0 24012 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_261
timestamp 1636968456
transform 1 0 25116 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_159_273
timestamp 1
transform 1 0 26220 0 -1 89216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_159_279
timestamp 1
transform 1 0 26772 0 -1 89216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_159_281
timestamp 1636968456
transform 1 0 26956 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_293
timestamp 1636968456
transform 1 0 28060 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_305
timestamp 1636968456
transform 1 0 29164 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_317
timestamp 1636968456
transform 1 0 30268 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_159_329
timestamp 1
transform 1 0 31372 0 -1 89216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_159_335
timestamp 1
transform 1 0 31924 0 -1 89216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_159_337
timestamp 1636968456
transform 1 0 32108 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_349
timestamp 1636968456
transform 1 0 33212 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_361
timestamp 1636968456
transform 1 0 34316 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_373
timestamp 1636968456
transform 1 0 35420 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_159_385
timestamp 1
transform 1 0 36524 0 -1 89216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_159_391
timestamp 1
transform 1 0 37076 0 -1 89216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_159_393
timestamp 1636968456
transform 1 0 37260 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_405
timestamp 1636968456
transform 1 0 38364 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_417
timestamp 1636968456
transform 1 0 39468 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_429
timestamp 1636968456
transform 1 0 40572 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_159_441
timestamp 1
transform 1 0 41676 0 -1 89216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_159_447
timestamp 1
transform 1 0 42228 0 -1 89216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_159_449
timestamp 1636968456
transform 1 0 42412 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_461
timestamp 1636968456
transform 1 0 43516 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_473
timestamp 1636968456
transform 1 0 44620 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_485
timestamp 1636968456
transform 1 0 45724 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_159_497
timestamp 1
transform 1 0 46828 0 -1 89216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_159_503
timestamp 1
transform 1 0 47380 0 -1 89216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_159_505
timestamp 1636968456
transform 1 0 47564 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_517
timestamp 1636968456
transform 1 0 48668 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_529
timestamp 1636968456
transform 1 0 49772 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_541
timestamp 1636968456
transform 1 0 50876 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_159_553
timestamp 1
transform 1 0 51980 0 -1 89216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_159_559
timestamp 1
transform 1 0 52532 0 -1 89216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_159_561
timestamp 1636968456
transform 1 0 52716 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_573
timestamp 1636968456
transform 1 0 53820 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_585
timestamp 1636968456
transform 1 0 54924 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_597
timestamp 1636968456
transform 1 0 56028 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_159_609
timestamp 1
transform 1 0 57132 0 -1 89216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_159_615
timestamp 1
transform 1 0 57684 0 -1 89216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_159_617
timestamp 1636968456
transform 1 0 57868 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_629
timestamp 1636968456
transform 1 0 58972 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_641
timestamp 1636968456
transform 1 0 60076 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_653
timestamp 1636968456
transform 1 0 61180 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_159_665
timestamp 1
transform 1 0 62284 0 -1 89216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_159_671
timestamp 1
transform 1 0 62836 0 -1 89216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_159_673
timestamp 1636968456
transform 1 0 63020 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_685
timestamp 1636968456
transform 1 0 64124 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_697
timestamp 1636968456
transform 1 0 65228 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_709
timestamp 1636968456
transform 1 0 66332 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_159_721
timestamp 1
transform 1 0 67436 0 -1 89216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_159_727
timestamp 1
transform 1 0 67988 0 -1 89216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_159_729
timestamp 1636968456
transform 1 0 68172 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_741
timestamp 1636968456
transform 1 0 69276 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_753
timestamp 1636968456
transform 1 0 70380 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_765
timestamp 1636968456
transform 1 0 71484 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_159_777
timestamp 1
transform 1 0 72588 0 -1 89216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_159_783
timestamp 1
transform 1 0 73140 0 -1 89216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_159_785
timestamp 1636968456
transform 1 0 73324 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_797
timestamp 1636968456
transform 1 0 74428 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_809
timestamp 1636968456
transform 1 0 75532 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_821
timestamp 1636968456
transform 1 0 76636 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_159_833
timestamp 1
transform 1 0 77740 0 -1 89216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_159_839
timestamp 1
transform 1 0 78292 0 -1 89216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_159_841
timestamp 1636968456
transform 1 0 78476 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_853
timestamp 1636968456
transform 1 0 79580 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_865
timestamp 1636968456
transform 1 0 80684 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_877
timestamp 1636968456
transform 1 0 81788 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_159_889
timestamp 1
transform 1 0 82892 0 -1 89216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_159_895
timestamp 1
transform 1 0 83444 0 -1 89216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_159_897
timestamp 1636968456
transform 1 0 83628 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_909
timestamp 1636968456
transform 1 0 84732 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_921
timestamp 1636968456
transform 1 0 85836 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_933
timestamp 1636968456
transform 1 0 86940 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_159_945
timestamp 1
transform 1 0 88044 0 -1 89216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_159_951
timestamp 1
transform 1 0 88596 0 -1 89216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_159_953
timestamp 1636968456
transform 1 0 88780 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_965
timestamp 1636968456
transform 1 0 89884 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_977
timestamp 1636968456
transform 1 0 90988 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_989
timestamp 1636968456
transform 1 0 92092 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_159_1001
timestamp 1
transform 1 0 93196 0 -1 89216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_159_1007
timestamp 1
transform 1 0 93748 0 -1 89216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_159_1009
timestamp 1636968456
transform 1 0 93932 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_1021
timestamp 1636968456
transform 1 0 95036 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_1033
timestamp 1636968456
transform 1 0 96140 0 -1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_159_1045
timestamp 1636968456
transform 1 0 97244 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_159_1057
timestamp 1
transform 1 0 98348 0 -1 89216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_159_1063
timestamp 1
transform 1 0 98900 0 -1 89216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_159_1065
timestamp 1636968456
transform 1 0 99084 0 -1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_159_1077
timestamp 1
transform 1 0 100188 0 -1 89216
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_160_3
timestamp 1636968456
transform 1 0 1380 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_15
timestamp 1636968456
transform 1 0 2484 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_160_27
timestamp 1
transform 1 0 3588 0 1 89216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_160_29
timestamp 1636968456
transform 1 0 3772 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_41
timestamp 1636968456
transform 1 0 4876 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_53
timestamp 1636968456
transform 1 0 5980 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_65
timestamp 1636968456
transform 1 0 7084 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_160_77
timestamp 1
transform 1 0 8188 0 1 89216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_160_83
timestamp 1
transform 1 0 8740 0 1 89216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_160_85
timestamp 1636968456
transform 1 0 8924 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_97
timestamp 1636968456
transform 1 0 10028 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_109
timestamp 1636968456
transform 1 0 11132 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_121
timestamp 1636968456
transform 1 0 12236 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_160_133
timestamp 1
transform 1 0 13340 0 1 89216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_160_139
timestamp 1
transform 1 0 13892 0 1 89216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_160_141
timestamp 1636968456
transform 1 0 14076 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_153
timestamp 1636968456
transform 1 0 15180 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_165
timestamp 1636968456
transform 1 0 16284 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_177
timestamp 1636968456
transform 1 0 17388 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_160_189
timestamp 1
transform 1 0 18492 0 1 89216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_160_195
timestamp 1
transform 1 0 19044 0 1 89216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_160_197
timestamp 1636968456
transform 1 0 19228 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_209
timestamp 1636968456
transform 1 0 20332 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_221
timestamp 1636968456
transform 1 0 21436 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_233
timestamp 1636968456
transform 1 0 22540 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_160_245
timestamp 1
transform 1 0 23644 0 1 89216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_160_251
timestamp 1
transform 1 0 24196 0 1 89216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_160_253
timestamp 1636968456
transform 1 0 24380 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_265
timestamp 1636968456
transform 1 0 25484 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_277
timestamp 1636968456
transform 1 0 26588 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_289
timestamp 1636968456
transform 1 0 27692 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_160_301
timestamp 1
transform 1 0 28796 0 1 89216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_160_307
timestamp 1
transform 1 0 29348 0 1 89216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_160_309
timestamp 1636968456
transform 1 0 29532 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_321
timestamp 1636968456
transform 1 0 30636 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_333
timestamp 1636968456
transform 1 0 31740 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_345
timestamp 1636968456
transform 1 0 32844 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_160_357
timestamp 1
transform 1 0 33948 0 1 89216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_160_363
timestamp 1
transform 1 0 34500 0 1 89216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_160_365
timestamp 1636968456
transform 1 0 34684 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_377
timestamp 1636968456
transform 1 0 35788 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_389
timestamp 1636968456
transform 1 0 36892 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_401
timestamp 1636968456
transform 1 0 37996 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_160_413
timestamp 1
transform 1 0 39100 0 1 89216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_160_419
timestamp 1
transform 1 0 39652 0 1 89216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_160_421
timestamp 1636968456
transform 1 0 39836 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_433
timestamp 1636968456
transform 1 0 40940 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_445
timestamp 1636968456
transform 1 0 42044 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_457
timestamp 1636968456
transform 1 0 43148 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_160_469
timestamp 1
transform 1 0 44252 0 1 89216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_160_475
timestamp 1
transform 1 0 44804 0 1 89216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_160_477
timestamp 1636968456
transform 1 0 44988 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_489
timestamp 1636968456
transform 1 0 46092 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_501
timestamp 1636968456
transform 1 0 47196 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_513
timestamp 1636968456
transform 1 0 48300 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_160_525
timestamp 1
transform 1 0 49404 0 1 89216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_160_531
timestamp 1
transform 1 0 49956 0 1 89216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_160_533
timestamp 1636968456
transform 1 0 50140 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_545
timestamp 1636968456
transform 1 0 51244 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_557
timestamp 1636968456
transform 1 0 52348 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_569
timestamp 1636968456
transform 1 0 53452 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_160_581
timestamp 1
transform 1 0 54556 0 1 89216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_160_587
timestamp 1
transform 1 0 55108 0 1 89216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_160_589
timestamp 1636968456
transform 1 0 55292 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_601
timestamp 1636968456
transform 1 0 56396 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_613
timestamp 1636968456
transform 1 0 57500 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_625
timestamp 1636968456
transform 1 0 58604 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_160_637
timestamp 1
transform 1 0 59708 0 1 89216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_160_643
timestamp 1
transform 1 0 60260 0 1 89216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_160_645
timestamp 1636968456
transform 1 0 60444 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_657
timestamp 1636968456
transform 1 0 61548 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_669
timestamp 1636968456
transform 1 0 62652 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_681
timestamp 1636968456
transform 1 0 63756 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_160_693
timestamp 1
transform 1 0 64860 0 1 89216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_160_699
timestamp 1
transform 1 0 65412 0 1 89216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_160_701
timestamp 1636968456
transform 1 0 65596 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_713
timestamp 1636968456
transform 1 0 66700 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_725
timestamp 1636968456
transform 1 0 67804 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_737
timestamp 1636968456
transform 1 0 68908 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_160_749
timestamp 1
transform 1 0 70012 0 1 89216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_160_755
timestamp 1
transform 1 0 70564 0 1 89216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_160_757
timestamp 1636968456
transform 1 0 70748 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_769
timestamp 1636968456
transform 1 0 71852 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_781
timestamp 1636968456
transform 1 0 72956 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_793
timestamp 1636968456
transform 1 0 74060 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_160_805
timestamp 1
transform 1 0 75164 0 1 89216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_160_811
timestamp 1
transform 1 0 75716 0 1 89216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_160_813
timestamp 1636968456
transform 1 0 75900 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_825
timestamp 1636968456
transform 1 0 77004 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_837
timestamp 1636968456
transform 1 0 78108 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_849
timestamp 1636968456
transform 1 0 79212 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_160_861
timestamp 1
transform 1 0 80316 0 1 89216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_160_867
timestamp 1
transform 1 0 80868 0 1 89216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_160_869
timestamp 1636968456
transform 1 0 81052 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_881
timestamp 1636968456
transform 1 0 82156 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_893
timestamp 1636968456
transform 1 0 83260 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_905
timestamp 1636968456
transform 1 0 84364 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_160_917
timestamp 1
transform 1 0 85468 0 1 89216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_160_923
timestamp 1
transform 1 0 86020 0 1 89216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_160_925
timestamp 1636968456
transform 1 0 86204 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_937
timestamp 1636968456
transform 1 0 87308 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_949
timestamp 1636968456
transform 1 0 88412 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_961
timestamp 1636968456
transform 1 0 89516 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_160_973
timestamp 1
transform 1 0 90620 0 1 89216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_160_979
timestamp 1
transform 1 0 91172 0 1 89216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_160_981
timestamp 1636968456
transform 1 0 91356 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_993
timestamp 1636968456
transform 1 0 92460 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_1005
timestamp 1636968456
transform 1 0 93564 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_1017
timestamp 1636968456
transform 1 0 94668 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_160_1029
timestamp 1
transform 1 0 95772 0 1 89216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_160_1035
timestamp 1
transform 1 0 96324 0 1 89216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_160_1037
timestamp 1636968456
transform 1 0 96508 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_1049
timestamp 1636968456
transform 1 0 97612 0 1 89216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_160_1061
timestamp 1636968456
transform 1 0 98716 0 1 89216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_160_1073
timestamp 1
transform 1 0 99820 0 1 89216
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_161_3
timestamp 1636968456
transform 1 0 1380 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_15
timestamp 1636968456
transform 1 0 2484 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_27
timestamp 1636968456
transform 1 0 3588 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_39
timestamp 1636968456
transform 1 0 4692 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_161_51
timestamp 1
transform 1 0 5796 0 -1 90304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_161_55
timestamp 1
transform 1 0 6164 0 -1 90304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_161_57
timestamp 1636968456
transform 1 0 6348 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_69
timestamp 1636968456
transform 1 0 7452 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_81
timestamp 1636968456
transform 1 0 8556 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_93
timestamp 1636968456
transform 1 0 9660 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_161_105
timestamp 1
transform 1 0 10764 0 -1 90304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_161_111
timestamp 1
transform 1 0 11316 0 -1 90304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_161_113
timestamp 1636968456
transform 1 0 11500 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_125
timestamp 1636968456
transform 1 0 12604 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_137
timestamp 1636968456
transform 1 0 13708 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_149
timestamp 1636968456
transform 1 0 14812 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_161_161
timestamp 1
transform 1 0 15916 0 -1 90304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_161_167
timestamp 1
transform 1 0 16468 0 -1 90304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_161_169
timestamp 1636968456
transform 1 0 16652 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_181
timestamp 1636968456
transform 1 0 17756 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_193
timestamp 1636968456
transform 1 0 18860 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_205
timestamp 1636968456
transform 1 0 19964 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_161_217
timestamp 1
transform 1 0 21068 0 -1 90304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_161_223
timestamp 1
transform 1 0 21620 0 -1 90304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_161_225
timestamp 1636968456
transform 1 0 21804 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_237
timestamp 1636968456
transform 1 0 22908 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_249
timestamp 1636968456
transform 1 0 24012 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_261
timestamp 1636968456
transform 1 0 25116 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_161_273
timestamp 1
transform 1 0 26220 0 -1 90304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_161_279
timestamp 1
transform 1 0 26772 0 -1 90304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_161_281
timestamp 1636968456
transform 1 0 26956 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_293
timestamp 1636968456
transform 1 0 28060 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_305
timestamp 1636968456
transform 1 0 29164 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_317
timestamp 1636968456
transform 1 0 30268 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_161_329
timestamp 1
transform 1 0 31372 0 -1 90304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_161_335
timestamp 1
transform 1 0 31924 0 -1 90304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_161_337
timestamp 1636968456
transform 1 0 32108 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_349
timestamp 1636968456
transform 1 0 33212 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_361
timestamp 1636968456
transform 1 0 34316 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_373
timestamp 1636968456
transform 1 0 35420 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_161_385
timestamp 1
transform 1 0 36524 0 -1 90304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_161_391
timestamp 1
transform 1 0 37076 0 -1 90304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_161_393
timestamp 1636968456
transform 1 0 37260 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_405
timestamp 1636968456
transform 1 0 38364 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_417
timestamp 1636968456
transform 1 0 39468 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_429
timestamp 1636968456
transform 1 0 40572 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_161_441
timestamp 1
transform 1 0 41676 0 -1 90304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_161_447
timestamp 1
transform 1 0 42228 0 -1 90304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_161_449
timestamp 1636968456
transform 1 0 42412 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_461
timestamp 1636968456
transform 1 0 43516 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_473
timestamp 1636968456
transform 1 0 44620 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_485
timestamp 1636968456
transform 1 0 45724 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_161_497
timestamp 1
transform 1 0 46828 0 -1 90304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_161_503
timestamp 1
transform 1 0 47380 0 -1 90304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_161_505
timestamp 1636968456
transform 1 0 47564 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_517
timestamp 1636968456
transform 1 0 48668 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_529
timestamp 1636968456
transform 1 0 49772 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_541
timestamp 1636968456
transform 1 0 50876 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_161_553
timestamp 1
transform 1 0 51980 0 -1 90304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_161_559
timestamp 1
transform 1 0 52532 0 -1 90304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_161_561
timestamp 1636968456
transform 1 0 52716 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_573
timestamp 1636968456
transform 1 0 53820 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_585
timestamp 1636968456
transform 1 0 54924 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_597
timestamp 1636968456
transform 1 0 56028 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_161_609
timestamp 1
transform 1 0 57132 0 -1 90304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_161_615
timestamp 1
transform 1 0 57684 0 -1 90304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_161_617
timestamp 1636968456
transform 1 0 57868 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_629
timestamp 1636968456
transform 1 0 58972 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_641
timestamp 1636968456
transform 1 0 60076 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_653
timestamp 1636968456
transform 1 0 61180 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_161_665
timestamp 1
transform 1 0 62284 0 -1 90304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_161_671
timestamp 1
transform 1 0 62836 0 -1 90304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_161_673
timestamp 1636968456
transform 1 0 63020 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_685
timestamp 1636968456
transform 1 0 64124 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_697
timestamp 1636968456
transform 1 0 65228 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_709
timestamp 1636968456
transform 1 0 66332 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_161_721
timestamp 1
transform 1 0 67436 0 -1 90304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_161_727
timestamp 1
transform 1 0 67988 0 -1 90304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_161_729
timestamp 1636968456
transform 1 0 68172 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_741
timestamp 1636968456
transform 1 0 69276 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_753
timestamp 1636968456
transform 1 0 70380 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_765
timestamp 1636968456
transform 1 0 71484 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_161_777
timestamp 1
transform 1 0 72588 0 -1 90304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_161_783
timestamp 1
transform 1 0 73140 0 -1 90304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_161_785
timestamp 1636968456
transform 1 0 73324 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_797
timestamp 1636968456
transform 1 0 74428 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_809
timestamp 1636968456
transform 1 0 75532 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_821
timestamp 1636968456
transform 1 0 76636 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_161_833
timestamp 1
transform 1 0 77740 0 -1 90304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_161_839
timestamp 1
transform 1 0 78292 0 -1 90304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_161_841
timestamp 1636968456
transform 1 0 78476 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_853
timestamp 1636968456
transform 1 0 79580 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_865
timestamp 1636968456
transform 1 0 80684 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_877
timestamp 1636968456
transform 1 0 81788 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_161_889
timestamp 1
transform 1 0 82892 0 -1 90304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_161_895
timestamp 1
transform 1 0 83444 0 -1 90304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_161_897
timestamp 1636968456
transform 1 0 83628 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_909
timestamp 1636968456
transform 1 0 84732 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_921
timestamp 1636968456
transform 1 0 85836 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_933
timestamp 1636968456
transform 1 0 86940 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_161_945
timestamp 1
transform 1 0 88044 0 -1 90304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_161_951
timestamp 1
transform 1 0 88596 0 -1 90304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_161_953
timestamp 1636968456
transform 1 0 88780 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_965
timestamp 1636968456
transform 1 0 89884 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_977
timestamp 1636968456
transform 1 0 90988 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_989
timestamp 1636968456
transform 1 0 92092 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_161_1001
timestamp 1
transform 1 0 93196 0 -1 90304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_161_1007
timestamp 1
transform 1 0 93748 0 -1 90304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_161_1009
timestamp 1636968456
transform 1 0 93932 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_1021
timestamp 1636968456
transform 1 0 95036 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_1033
timestamp 1636968456
transform 1 0 96140 0 -1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_161_1045
timestamp 1636968456
transform 1 0 97244 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_161_1057
timestamp 1
transform 1 0 98348 0 -1 90304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_161_1063
timestamp 1
transform 1 0 98900 0 -1 90304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_161_1065
timestamp 1636968456
transform 1 0 99084 0 -1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_161_1077
timestamp 1
transform 1 0 100188 0 -1 90304
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_162_3
timestamp 1636968456
transform 1 0 1380 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_15
timestamp 1636968456
transform 1 0 2484 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_162_27
timestamp 1
transform 1 0 3588 0 1 90304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_162_29
timestamp 1636968456
transform 1 0 3772 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_41
timestamp 1636968456
transform 1 0 4876 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_53
timestamp 1636968456
transform 1 0 5980 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_65
timestamp 1636968456
transform 1 0 7084 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_162_77
timestamp 1
transform 1 0 8188 0 1 90304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_162_83
timestamp 1
transform 1 0 8740 0 1 90304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_162_85
timestamp 1636968456
transform 1 0 8924 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_97
timestamp 1636968456
transform 1 0 10028 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_109
timestamp 1636968456
transform 1 0 11132 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_121
timestamp 1636968456
transform 1 0 12236 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_162_133
timestamp 1
transform 1 0 13340 0 1 90304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_162_139
timestamp 1
transform 1 0 13892 0 1 90304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_162_141
timestamp 1636968456
transform 1 0 14076 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_153
timestamp 1636968456
transform 1 0 15180 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_165
timestamp 1636968456
transform 1 0 16284 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_177
timestamp 1636968456
transform 1 0 17388 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_162_189
timestamp 1
transform 1 0 18492 0 1 90304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_162_195
timestamp 1
transform 1 0 19044 0 1 90304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_162_197
timestamp 1636968456
transform 1 0 19228 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_209
timestamp 1636968456
transform 1 0 20332 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_221
timestamp 1636968456
transform 1 0 21436 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_233
timestamp 1636968456
transform 1 0 22540 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_162_245
timestamp 1
transform 1 0 23644 0 1 90304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_162_251
timestamp 1
transform 1 0 24196 0 1 90304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_162_253
timestamp 1636968456
transform 1 0 24380 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_265
timestamp 1636968456
transform 1 0 25484 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_277
timestamp 1636968456
transform 1 0 26588 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_289
timestamp 1636968456
transform 1 0 27692 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_162_301
timestamp 1
transform 1 0 28796 0 1 90304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_162_307
timestamp 1
transform 1 0 29348 0 1 90304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_162_309
timestamp 1636968456
transform 1 0 29532 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_321
timestamp 1636968456
transform 1 0 30636 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_333
timestamp 1636968456
transform 1 0 31740 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_345
timestamp 1636968456
transform 1 0 32844 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_162_357
timestamp 1
transform 1 0 33948 0 1 90304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_162_363
timestamp 1
transform 1 0 34500 0 1 90304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_162_365
timestamp 1636968456
transform 1 0 34684 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_377
timestamp 1636968456
transform 1 0 35788 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_389
timestamp 1636968456
transform 1 0 36892 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_401
timestamp 1636968456
transform 1 0 37996 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_162_413
timestamp 1
transform 1 0 39100 0 1 90304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_162_419
timestamp 1
transform 1 0 39652 0 1 90304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_162_421
timestamp 1636968456
transform 1 0 39836 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_433
timestamp 1636968456
transform 1 0 40940 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_445
timestamp 1636968456
transform 1 0 42044 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_457
timestamp 1636968456
transform 1 0 43148 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_162_469
timestamp 1
transform 1 0 44252 0 1 90304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_162_475
timestamp 1
transform 1 0 44804 0 1 90304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_162_477
timestamp 1636968456
transform 1 0 44988 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_489
timestamp 1636968456
transform 1 0 46092 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_501
timestamp 1636968456
transform 1 0 47196 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_513
timestamp 1636968456
transform 1 0 48300 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_162_525
timestamp 1
transform 1 0 49404 0 1 90304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_162_531
timestamp 1
transform 1 0 49956 0 1 90304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_162_533
timestamp 1636968456
transform 1 0 50140 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_545
timestamp 1636968456
transform 1 0 51244 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_557
timestamp 1636968456
transform 1 0 52348 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_569
timestamp 1636968456
transform 1 0 53452 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_162_581
timestamp 1
transform 1 0 54556 0 1 90304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_162_587
timestamp 1
transform 1 0 55108 0 1 90304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_162_589
timestamp 1636968456
transform 1 0 55292 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_601
timestamp 1636968456
transform 1 0 56396 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_613
timestamp 1636968456
transform 1 0 57500 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_625
timestamp 1636968456
transform 1 0 58604 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_162_637
timestamp 1
transform 1 0 59708 0 1 90304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_162_643
timestamp 1
transform 1 0 60260 0 1 90304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_162_645
timestamp 1636968456
transform 1 0 60444 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_657
timestamp 1636968456
transform 1 0 61548 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_669
timestamp 1636968456
transform 1 0 62652 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_681
timestamp 1636968456
transform 1 0 63756 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_162_693
timestamp 1
transform 1 0 64860 0 1 90304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_162_699
timestamp 1
transform 1 0 65412 0 1 90304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_162_701
timestamp 1636968456
transform 1 0 65596 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_713
timestamp 1636968456
transform 1 0 66700 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_725
timestamp 1636968456
transform 1 0 67804 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_737
timestamp 1636968456
transform 1 0 68908 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_162_749
timestamp 1
transform 1 0 70012 0 1 90304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_162_755
timestamp 1
transform 1 0 70564 0 1 90304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_162_757
timestamp 1636968456
transform 1 0 70748 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_769
timestamp 1636968456
transform 1 0 71852 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_781
timestamp 1636968456
transform 1 0 72956 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_793
timestamp 1636968456
transform 1 0 74060 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_162_805
timestamp 1
transform 1 0 75164 0 1 90304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_162_811
timestamp 1
transform 1 0 75716 0 1 90304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_162_813
timestamp 1636968456
transform 1 0 75900 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_825
timestamp 1636968456
transform 1 0 77004 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_837
timestamp 1636968456
transform 1 0 78108 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_849
timestamp 1636968456
transform 1 0 79212 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_162_861
timestamp 1
transform 1 0 80316 0 1 90304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_162_867
timestamp 1
transform 1 0 80868 0 1 90304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_162_869
timestamp 1636968456
transform 1 0 81052 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_881
timestamp 1636968456
transform 1 0 82156 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_893
timestamp 1636968456
transform 1 0 83260 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_905
timestamp 1636968456
transform 1 0 84364 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_162_917
timestamp 1
transform 1 0 85468 0 1 90304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_162_923
timestamp 1
transform 1 0 86020 0 1 90304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_162_925
timestamp 1636968456
transform 1 0 86204 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_937
timestamp 1636968456
transform 1 0 87308 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_949
timestamp 1636968456
transform 1 0 88412 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_961
timestamp 1636968456
transform 1 0 89516 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_162_973
timestamp 1
transform 1 0 90620 0 1 90304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_162_979
timestamp 1
transform 1 0 91172 0 1 90304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_162_981
timestamp 1636968456
transform 1 0 91356 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_993
timestamp 1636968456
transform 1 0 92460 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_1005
timestamp 1636968456
transform 1 0 93564 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_1017
timestamp 1636968456
transform 1 0 94668 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_162_1029
timestamp 1
transform 1 0 95772 0 1 90304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_162_1035
timestamp 1
transform 1 0 96324 0 1 90304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_162_1037
timestamp 1636968456
transform 1 0 96508 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_1049
timestamp 1636968456
transform 1 0 97612 0 1 90304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_162_1061
timestamp 1636968456
transform 1 0 98716 0 1 90304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_162_1073
timestamp 1
transform 1 0 99820 0 1 90304
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_163_3
timestamp 1636968456
transform 1 0 1380 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_15
timestamp 1636968456
transform 1 0 2484 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_27
timestamp 1636968456
transform 1 0 3588 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_39
timestamp 1636968456
transform 1 0 4692 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_163_51
timestamp 1
transform 1 0 5796 0 -1 91392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_163_55
timestamp 1
transform 1 0 6164 0 -1 91392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_163_57
timestamp 1636968456
transform 1 0 6348 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_69
timestamp 1636968456
transform 1 0 7452 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_81
timestamp 1636968456
transform 1 0 8556 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_93
timestamp 1636968456
transform 1 0 9660 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_163_105
timestamp 1
transform 1 0 10764 0 -1 91392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_163_111
timestamp 1
transform 1 0 11316 0 -1 91392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_163_113
timestamp 1636968456
transform 1 0 11500 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_125
timestamp 1636968456
transform 1 0 12604 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_137
timestamp 1636968456
transform 1 0 13708 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_149
timestamp 1636968456
transform 1 0 14812 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_163_161
timestamp 1
transform 1 0 15916 0 -1 91392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_163_167
timestamp 1
transform 1 0 16468 0 -1 91392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_163_169
timestamp 1636968456
transform 1 0 16652 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_181
timestamp 1636968456
transform 1 0 17756 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_193
timestamp 1636968456
transform 1 0 18860 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_205
timestamp 1636968456
transform 1 0 19964 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_163_217
timestamp 1
transform 1 0 21068 0 -1 91392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_163_223
timestamp 1
transform 1 0 21620 0 -1 91392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_163_225
timestamp 1636968456
transform 1 0 21804 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_237
timestamp 1636968456
transform 1 0 22908 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_249
timestamp 1636968456
transform 1 0 24012 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_261
timestamp 1636968456
transform 1 0 25116 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_163_273
timestamp 1
transform 1 0 26220 0 -1 91392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_163_279
timestamp 1
transform 1 0 26772 0 -1 91392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_163_281
timestamp 1636968456
transform 1 0 26956 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_293
timestamp 1636968456
transform 1 0 28060 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_305
timestamp 1636968456
transform 1 0 29164 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_317
timestamp 1636968456
transform 1 0 30268 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_163_329
timestamp 1
transform 1 0 31372 0 -1 91392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_163_335
timestamp 1
transform 1 0 31924 0 -1 91392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_163_337
timestamp 1636968456
transform 1 0 32108 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_349
timestamp 1636968456
transform 1 0 33212 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_361
timestamp 1636968456
transform 1 0 34316 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_373
timestamp 1636968456
transform 1 0 35420 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_163_385
timestamp 1
transform 1 0 36524 0 -1 91392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_163_391
timestamp 1
transform 1 0 37076 0 -1 91392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_163_393
timestamp 1636968456
transform 1 0 37260 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_405
timestamp 1636968456
transform 1 0 38364 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_417
timestamp 1636968456
transform 1 0 39468 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_429
timestamp 1636968456
transform 1 0 40572 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_163_441
timestamp 1
transform 1 0 41676 0 -1 91392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_163_447
timestamp 1
transform 1 0 42228 0 -1 91392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_163_449
timestamp 1636968456
transform 1 0 42412 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_461
timestamp 1636968456
transform 1 0 43516 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_473
timestamp 1636968456
transform 1 0 44620 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_485
timestamp 1636968456
transform 1 0 45724 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_163_497
timestamp 1
transform 1 0 46828 0 -1 91392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_163_503
timestamp 1
transform 1 0 47380 0 -1 91392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_163_505
timestamp 1636968456
transform 1 0 47564 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_517
timestamp 1636968456
transform 1 0 48668 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_529
timestamp 1636968456
transform 1 0 49772 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_541
timestamp 1636968456
transform 1 0 50876 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_163_553
timestamp 1
transform 1 0 51980 0 -1 91392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_163_559
timestamp 1
transform 1 0 52532 0 -1 91392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_163_561
timestamp 1636968456
transform 1 0 52716 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_573
timestamp 1636968456
transform 1 0 53820 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_585
timestamp 1636968456
transform 1 0 54924 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_597
timestamp 1636968456
transform 1 0 56028 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_163_609
timestamp 1
transform 1 0 57132 0 -1 91392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_163_615
timestamp 1
transform 1 0 57684 0 -1 91392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_163_617
timestamp 1636968456
transform 1 0 57868 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_629
timestamp 1636968456
transform 1 0 58972 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_641
timestamp 1636968456
transform 1 0 60076 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_653
timestamp 1636968456
transform 1 0 61180 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_163_665
timestamp 1
transform 1 0 62284 0 -1 91392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_163_671
timestamp 1
transform 1 0 62836 0 -1 91392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_163_673
timestamp 1636968456
transform 1 0 63020 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_685
timestamp 1636968456
transform 1 0 64124 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_697
timestamp 1636968456
transform 1 0 65228 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_709
timestamp 1636968456
transform 1 0 66332 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_163_721
timestamp 1
transform 1 0 67436 0 -1 91392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_163_727
timestamp 1
transform 1 0 67988 0 -1 91392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_163_729
timestamp 1636968456
transform 1 0 68172 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_741
timestamp 1636968456
transform 1 0 69276 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_753
timestamp 1636968456
transform 1 0 70380 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_765
timestamp 1636968456
transform 1 0 71484 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_163_777
timestamp 1
transform 1 0 72588 0 -1 91392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_163_783
timestamp 1
transform 1 0 73140 0 -1 91392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_163_785
timestamp 1636968456
transform 1 0 73324 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_797
timestamp 1636968456
transform 1 0 74428 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_809
timestamp 1636968456
transform 1 0 75532 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_821
timestamp 1636968456
transform 1 0 76636 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_163_833
timestamp 1
transform 1 0 77740 0 -1 91392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_163_839
timestamp 1
transform 1 0 78292 0 -1 91392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_163_841
timestamp 1636968456
transform 1 0 78476 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_853
timestamp 1636968456
transform 1 0 79580 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_865
timestamp 1636968456
transform 1 0 80684 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_877
timestamp 1636968456
transform 1 0 81788 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_163_889
timestamp 1
transform 1 0 82892 0 -1 91392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_163_895
timestamp 1
transform 1 0 83444 0 -1 91392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_163_897
timestamp 1636968456
transform 1 0 83628 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_909
timestamp 1636968456
transform 1 0 84732 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_921
timestamp 1636968456
transform 1 0 85836 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_933
timestamp 1636968456
transform 1 0 86940 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_163_945
timestamp 1
transform 1 0 88044 0 -1 91392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_163_951
timestamp 1
transform 1 0 88596 0 -1 91392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_163_953
timestamp 1636968456
transform 1 0 88780 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_965
timestamp 1636968456
transform 1 0 89884 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_977
timestamp 1636968456
transform 1 0 90988 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_989
timestamp 1636968456
transform 1 0 92092 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_163_1001
timestamp 1
transform 1 0 93196 0 -1 91392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_163_1007
timestamp 1
transform 1 0 93748 0 -1 91392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_163_1009
timestamp 1636968456
transform 1 0 93932 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_1021
timestamp 1636968456
transform 1 0 95036 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_1033
timestamp 1636968456
transform 1 0 96140 0 -1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_163_1045
timestamp 1636968456
transform 1 0 97244 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_163_1057
timestamp 1
transform 1 0 98348 0 -1 91392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_163_1063
timestamp 1
transform 1 0 98900 0 -1 91392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_163_1065
timestamp 1636968456
transform 1 0 99084 0 -1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_163_1077
timestamp 1
transform 1 0 100188 0 -1 91392
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_164_3
timestamp 1636968456
transform 1 0 1380 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_15
timestamp 1636968456
transform 1 0 2484 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_164_27
timestamp 1
transform 1 0 3588 0 1 91392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_164_29
timestamp 1636968456
transform 1 0 3772 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_41
timestamp 1636968456
transform 1 0 4876 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_53
timestamp 1636968456
transform 1 0 5980 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_65
timestamp 1636968456
transform 1 0 7084 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_164_77
timestamp 1
transform 1 0 8188 0 1 91392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_164_83
timestamp 1
transform 1 0 8740 0 1 91392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_164_85
timestamp 1636968456
transform 1 0 8924 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_97
timestamp 1636968456
transform 1 0 10028 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_109
timestamp 1636968456
transform 1 0 11132 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_121
timestamp 1636968456
transform 1 0 12236 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_164_133
timestamp 1
transform 1 0 13340 0 1 91392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_164_139
timestamp 1
transform 1 0 13892 0 1 91392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_164_141
timestamp 1636968456
transform 1 0 14076 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_153
timestamp 1636968456
transform 1 0 15180 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_165
timestamp 1636968456
transform 1 0 16284 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_177
timestamp 1636968456
transform 1 0 17388 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_164_189
timestamp 1
transform 1 0 18492 0 1 91392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_164_195
timestamp 1
transform 1 0 19044 0 1 91392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_164_197
timestamp 1636968456
transform 1 0 19228 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_209
timestamp 1636968456
transform 1 0 20332 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_221
timestamp 1636968456
transform 1 0 21436 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_233
timestamp 1636968456
transform 1 0 22540 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_164_245
timestamp 1
transform 1 0 23644 0 1 91392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_164_251
timestamp 1
transform 1 0 24196 0 1 91392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_164_253
timestamp 1636968456
transform 1 0 24380 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_265
timestamp 1636968456
transform 1 0 25484 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_277
timestamp 1636968456
transform 1 0 26588 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_289
timestamp 1636968456
transform 1 0 27692 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_164_301
timestamp 1
transform 1 0 28796 0 1 91392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_164_307
timestamp 1
transform 1 0 29348 0 1 91392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_164_309
timestamp 1636968456
transform 1 0 29532 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_321
timestamp 1636968456
transform 1 0 30636 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_333
timestamp 1636968456
transform 1 0 31740 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_345
timestamp 1636968456
transform 1 0 32844 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_164_357
timestamp 1
transform 1 0 33948 0 1 91392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_164_363
timestamp 1
transform 1 0 34500 0 1 91392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_164_365
timestamp 1636968456
transform 1 0 34684 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_377
timestamp 1636968456
transform 1 0 35788 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_389
timestamp 1636968456
transform 1 0 36892 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_401
timestamp 1636968456
transform 1 0 37996 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_164_413
timestamp 1
transform 1 0 39100 0 1 91392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_164_419
timestamp 1
transform 1 0 39652 0 1 91392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_164_421
timestamp 1636968456
transform 1 0 39836 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_433
timestamp 1636968456
transform 1 0 40940 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_445
timestamp 1636968456
transform 1 0 42044 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_457
timestamp 1636968456
transform 1 0 43148 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_164_469
timestamp 1
transform 1 0 44252 0 1 91392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_164_475
timestamp 1
transform 1 0 44804 0 1 91392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_164_477
timestamp 1636968456
transform 1 0 44988 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_489
timestamp 1636968456
transform 1 0 46092 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_501
timestamp 1636968456
transform 1 0 47196 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_513
timestamp 1636968456
transform 1 0 48300 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_164_525
timestamp 1
transform 1 0 49404 0 1 91392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_164_531
timestamp 1
transform 1 0 49956 0 1 91392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_164_533
timestamp 1636968456
transform 1 0 50140 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_545
timestamp 1636968456
transform 1 0 51244 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_557
timestamp 1636968456
transform 1 0 52348 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_569
timestamp 1636968456
transform 1 0 53452 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_164_581
timestamp 1
transform 1 0 54556 0 1 91392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_164_587
timestamp 1
transform 1 0 55108 0 1 91392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_164_589
timestamp 1636968456
transform 1 0 55292 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_601
timestamp 1636968456
transform 1 0 56396 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_613
timestamp 1636968456
transform 1 0 57500 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_625
timestamp 1636968456
transform 1 0 58604 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_164_637
timestamp 1
transform 1 0 59708 0 1 91392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_164_643
timestamp 1
transform 1 0 60260 0 1 91392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_164_645
timestamp 1636968456
transform 1 0 60444 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_657
timestamp 1636968456
transform 1 0 61548 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_669
timestamp 1636968456
transform 1 0 62652 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_681
timestamp 1636968456
transform 1 0 63756 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_164_693
timestamp 1
transform 1 0 64860 0 1 91392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_164_699
timestamp 1
transform 1 0 65412 0 1 91392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_164_701
timestamp 1636968456
transform 1 0 65596 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_713
timestamp 1636968456
transform 1 0 66700 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_725
timestamp 1636968456
transform 1 0 67804 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_737
timestamp 1636968456
transform 1 0 68908 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_164_749
timestamp 1
transform 1 0 70012 0 1 91392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_164_755
timestamp 1
transform 1 0 70564 0 1 91392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_164_757
timestamp 1636968456
transform 1 0 70748 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_769
timestamp 1636968456
transform 1 0 71852 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_781
timestamp 1636968456
transform 1 0 72956 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_793
timestamp 1636968456
transform 1 0 74060 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_164_805
timestamp 1
transform 1 0 75164 0 1 91392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_164_811
timestamp 1
transform 1 0 75716 0 1 91392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_164_813
timestamp 1636968456
transform 1 0 75900 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_825
timestamp 1636968456
transform 1 0 77004 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_837
timestamp 1636968456
transform 1 0 78108 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_849
timestamp 1636968456
transform 1 0 79212 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_164_861
timestamp 1
transform 1 0 80316 0 1 91392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_164_867
timestamp 1
transform 1 0 80868 0 1 91392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_164_869
timestamp 1636968456
transform 1 0 81052 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_881
timestamp 1636968456
transform 1 0 82156 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_893
timestamp 1636968456
transform 1 0 83260 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_905
timestamp 1636968456
transform 1 0 84364 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_164_917
timestamp 1
transform 1 0 85468 0 1 91392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_164_923
timestamp 1
transform 1 0 86020 0 1 91392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_164_925
timestamp 1636968456
transform 1 0 86204 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_937
timestamp 1636968456
transform 1 0 87308 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_949
timestamp 1636968456
transform 1 0 88412 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_961
timestamp 1636968456
transform 1 0 89516 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_164_973
timestamp 1
transform 1 0 90620 0 1 91392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_164_979
timestamp 1
transform 1 0 91172 0 1 91392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_164_981
timestamp 1636968456
transform 1 0 91356 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_993
timestamp 1636968456
transform 1 0 92460 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_1005
timestamp 1636968456
transform 1 0 93564 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_1017
timestamp 1636968456
transform 1 0 94668 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_164_1029
timestamp 1
transform 1 0 95772 0 1 91392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_164_1035
timestamp 1
transform 1 0 96324 0 1 91392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_164_1037
timestamp 1636968456
transform 1 0 96508 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_1049
timestamp 1636968456
transform 1 0 97612 0 1 91392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_164_1061
timestamp 1636968456
transform 1 0 98716 0 1 91392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_164_1073
timestamp 1
transform 1 0 99820 0 1 91392
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_165_3
timestamp 1636968456
transform 1 0 1380 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_15
timestamp 1636968456
transform 1 0 2484 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_27
timestamp 1636968456
transform 1 0 3588 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_39
timestamp 1636968456
transform 1 0 4692 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_165_51
timestamp 1
transform 1 0 5796 0 -1 92480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_165_55
timestamp 1
transform 1 0 6164 0 -1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_165_57
timestamp 1636968456
transform 1 0 6348 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_69
timestamp 1636968456
transform 1 0 7452 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_81
timestamp 1636968456
transform 1 0 8556 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_93
timestamp 1636968456
transform 1 0 9660 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_165_105
timestamp 1
transform 1 0 10764 0 -1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_165_111
timestamp 1
transform 1 0 11316 0 -1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_165_113
timestamp 1636968456
transform 1 0 11500 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_125
timestamp 1636968456
transform 1 0 12604 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_137
timestamp 1636968456
transform 1 0 13708 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_149
timestamp 1636968456
transform 1 0 14812 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_165_161
timestamp 1
transform 1 0 15916 0 -1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_165_167
timestamp 1
transform 1 0 16468 0 -1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_165_169
timestamp 1636968456
transform 1 0 16652 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_181
timestamp 1636968456
transform 1 0 17756 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_193
timestamp 1636968456
transform 1 0 18860 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_205
timestamp 1636968456
transform 1 0 19964 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_165_217
timestamp 1
transform 1 0 21068 0 -1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_165_223
timestamp 1
transform 1 0 21620 0 -1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_165_225
timestamp 1636968456
transform 1 0 21804 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_237
timestamp 1636968456
transform 1 0 22908 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_249
timestamp 1636968456
transform 1 0 24012 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_261
timestamp 1636968456
transform 1 0 25116 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_165_273
timestamp 1
transform 1 0 26220 0 -1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_165_279
timestamp 1
transform 1 0 26772 0 -1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_165_281
timestamp 1636968456
transform 1 0 26956 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_293
timestamp 1636968456
transform 1 0 28060 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_305
timestamp 1636968456
transform 1 0 29164 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_317
timestamp 1636968456
transform 1 0 30268 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_165_329
timestamp 1
transform 1 0 31372 0 -1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_165_335
timestamp 1
transform 1 0 31924 0 -1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_165_337
timestamp 1636968456
transform 1 0 32108 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_349
timestamp 1636968456
transform 1 0 33212 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_361
timestamp 1636968456
transform 1 0 34316 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_373
timestamp 1636968456
transform 1 0 35420 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_165_385
timestamp 1
transform 1 0 36524 0 -1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_165_391
timestamp 1
transform 1 0 37076 0 -1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_165_393
timestamp 1636968456
transform 1 0 37260 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_405
timestamp 1636968456
transform 1 0 38364 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_417
timestamp 1636968456
transform 1 0 39468 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_429
timestamp 1636968456
transform 1 0 40572 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_165_441
timestamp 1
transform 1 0 41676 0 -1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_165_447
timestamp 1
transform 1 0 42228 0 -1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_165_449
timestamp 1636968456
transform 1 0 42412 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_461
timestamp 1636968456
transform 1 0 43516 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_473
timestamp 1636968456
transform 1 0 44620 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_485
timestamp 1636968456
transform 1 0 45724 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_165_497
timestamp 1
transform 1 0 46828 0 -1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_165_503
timestamp 1
transform 1 0 47380 0 -1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_165_505
timestamp 1636968456
transform 1 0 47564 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_517
timestamp 1636968456
transform 1 0 48668 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_529
timestamp 1636968456
transform 1 0 49772 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_541
timestamp 1636968456
transform 1 0 50876 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_165_553
timestamp 1
transform 1 0 51980 0 -1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_165_559
timestamp 1
transform 1 0 52532 0 -1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_165_561
timestamp 1636968456
transform 1 0 52716 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_573
timestamp 1636968456
transform 1 0 53820 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_585
timestamp 1636968456
transform 1 0 54924 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_597
timestamp 1636968456
transform 1 0 56028 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_165_609
timestamp 1
transform 1 0 57132 0 -1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_165_615
timestamp 1
transform 1 0 57684 0 -1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_165_617
timestamp 1636968456
transform 1 0 57868 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_629
timestamp 1636968456
transform 1 0 58972 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_641
timestamp 1636968456
transform 1 0 60076 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_653
timestamp 1636968456
transform 1 0 61180 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_165_665
timestamp 1
transform 1 0 62284 0 -1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_165_671
timestamp 1
transform 1 0 62836 0 -1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_165_673
timestamp 1636968456
transform 1 0 63020 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_685
timestamp 1636968456
transform 1 0 64124 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_697
timestamp 1636968456
transform 1 0 65228 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_709
timestamp 1636968456
transform 1 0 66332 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_165_721
timestamp 1
transform 1 0 67436 0 -1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_165_727
timestamp 1
transform 1 0 67988 0 -1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_165_729
timestamp 1636968456
transform 1 0 68172 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_741
timestamp 1636968456
transform 1 0 69276 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_753
timestamp 1636968456
transform 1 0 70380 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_765
timestamp 1636968456
transform 1 0 71484 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_165_777
timestamp 1
transform 1 0 72588 0 -1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_165_783
timestamp 1
transform 1 0 73140 0 -1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_165_785
timestamp 1636968456
transform 1 0 73324 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_797
timestamp 1636968456
transform 1 0 74428 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_809
timestamp 1636968456
transform 1 0 75532 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_821
timestamp 1636968456
transform 1 0 76636 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_165_833
timestamp 1
transform 1 0 77740 0 -1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_165_839
timestamp 1
transform 1 0 78292 0 -1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_165_841
timestamp 1636968456
transform 1 0 78476 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_853
timestamp 1636968456
transform 1 0 79580 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_865
timestamp 1636968456
transform 1 0 80684 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_877
timestamp 1636968456
transform 1 0 81788 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_165_889
timestamp 1
transform 1 0 82892 0 -1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_165_895
timestamp 1
transform 1 0 83444 0 -1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_165_897
timestamp 1636968456
transform 1 0 83628 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_909
timestamp 1636968456
transform 1 0 84732 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_921
timestamp 1636968456
transform 1 0 85836 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_933
timestamp 1636968456
transform 1 0 86940 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_165_945
timestamp 1
transform 1 0 88044 0 -1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_165_951
timestamp 1
transform 1 0 88596 0 -1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_165_953
timestamp 1636968456
transform 1 0 88780 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_965
timestamp 1636968456
transform 1 0 89884 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_977
timestamp 1636968456
transform 1 0 90988 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_989
timestamp 1636968456
transform 1 0 92092 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_165_1001
timestamp 1
transform 1 0 93196 0 -1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_165_1007
timestamp 1
transform 1 0 93748 0 -1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_165_1009
timestamp 1636968456
transform 1 0 93932 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_1021
timestamp 1636968456
transform 1 0 95036 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_1033
timestamp 1636968456
transform 1 0 96140 0 -1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_165_1045
timestamp 1636968456
transform 1 0 97244 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_165_1057
timestamp 1
transform 1 0 98348 0 -1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_165_1063
timestamp 1
transform 1 0 98900 0 -1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_165_1065
timestamp 1636968456
transform 1 0 99084 0 -1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_165_1077
timestamp 1
transform 1 0 100188 0 -1 92480
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_166_3
timestamp 1636968456
transform 1 0 1380 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_15
timestamp 1636968456
transform 1 0 2484 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_166_27
timestamp 1
transform 1 0 3588 0 1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_166_29
timestamp 1636968456
transform 1 0 3772 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_41
timestamp 1636968456
transform 1 0 4876 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_53
timestamp 1636968456
transform 1 0 5980 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_65
timestamp 1636968456
transform 1 0 7084 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_77
timestamp 1
transform 1 0 8188 0 1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_83
timestamp 1
transform 1 0 8740 0 1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_166_85
timestamp 1636968456
transform 1 0 8924 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_97
timestamp 1636968456
transform 1 0 10028 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_109
timestamp 1636968456
transform 1 0 11132 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_121
timestamp 1636968456
transform 1 0 12236 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_133
timestamp 1
transform 1 0 13340 0 1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_139
timestamp 1
transform 1 0 13892 0 1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_166_141
timestamp 1636968456
transform 1 0 14076 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_153
timestamp 1636968456
transform 1 0 15180 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_165
timestamp 1636968456
transform 1 0 16284 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_177
timestamp 1636968456
transform 1 0 17388 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_189
timestamp 1
transform 1 0 18492 0 1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_195
timestamp 1
transform 1 0 19044 0 1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_166_197
timestamp 1636968456
transform 1 0 19228 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_209
timestamp 1636968456
transform 1 0 20332 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_221
timestamp 1636968456
transform 1 0 21436 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_233
timestamp 1636968456
transform 1 0 22540 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_245
timestamp 1
transform 1 0 23644 0 1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_251
timestamp 1
transform 1 0 24196 0 1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_166_253
timestamp 1636968456
transform 1 0 24380 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_265
timestamp 1636968456
transform 1 0 25484 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_277
timestamp 1636968456
transform 1 0 26588 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_289
timestamp 1636968456
transform 1 0 27692 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_301
timestamp 1
transform 1 0 28796 0 1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_307
timestamp 1
transform 1 0 29348 0 1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_166_309
timestamp 1636968456
transform 1 0 29532 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_321
timestamp 1636968456
transform 1 0 30636 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_333
timestamp 1636968456
transform 1 0 31740 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_345
timestamp 1636968456
transform 1 0 32844 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_357
timestamp 1
transform 1 0 33948 0 1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_363
timestamp 1
transform 1 0 34500 0 1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_166_365
timestamp 1636968456
transform 1 0 34684 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_377
timestamp 1636968456
transform 1 0 35788 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_389
timestamp 1636968456
transform 1 0 36892 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_401
timestamp 1636968456
transform 1 0 37996 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_413
timestamp 1
transform 1 0 39100 0 1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_419
timestamp 1
transform 1 0 39652 0 1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_166_421
timestamp 1636968456
transform 1 0 39836 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_433
timestamp 1636968456
transform 1 0 40940 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_445
timestamp 1636968456
transform 1 0 42044 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_457
timestamp 1636968456
transform 1 0 43148 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_469
timestamp 1
transform 1 0 44252 0 1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_475
timestamp 1
transform 1 0 44804 0 1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_166_477
timestamp 1636968456
transform 1 0 44988 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_489
timestamp 1636968456
transform 1 0 46092 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_501
timestamp 1636968456
transform 1 0 47196 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_513
timestamp 1636968456
transform 1 0 48300 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_525
timestamp 1
transform 1 0 49404 0 1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_531
timestamp 1
transform 1 0 49956 0 1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_166_533
timestamp 1636968456
transform 1 0 50140 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_545
timestamp 1636968456
transform 1 0 51244 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_557
timestamp 1636968456
transform 1 0 52348 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_569
timestamp 1636968456
transform 1 0 53452 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_581
timestamp 1
transform 1 0 54556 0 1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_587
timestamp 1
transform 1 0 55108 0 1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_166_589
timestamp 1636968456
transform 1 0 55292 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_601
timestamp 1636968456
transform 1 0 56396 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_613
timestamp 1636968456
transform 1 0 57500 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_625
timestamp 1636968456
transform 1 0 58604 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_637
timestamp 1
transform 1 0 59708 0 1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_643
timestamp 1
transform 1 0 60260 0 1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_166_645
timestamp 1636968456
transform 1 0 60444 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_657
timestamp 1636968456
transform 1 0 61548 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_669
timestamp 1636968456
transform 1 0 62652 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_681
timestamp 1636968456
transform 1 0 63756 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_693
timestamp 1
transform 1 0 64860 0 1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_699
timestamp 1
transform 1 0 65412 0 1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_166_701
timestamp 1636968456
transform 1 0 65596 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_713
timestamp 1636968456
transform 1 0 66700 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_725
timestamp 1636968456
transform 1 0 67804 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_737
timestamp 1636968456
transform 1 0 68908 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_749
timestamp 1
transform 1 0 70012 0 1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_755
timestamp 1
transform 1 0 70564 0 1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_166_757
timestamp 1636968456
transform 1 0 70748 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_769
timestamp 1636968456
transform 1 0 71852 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_781
timestamp 1636968456
transform 1 0 72956 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_793
timestamp 1636968456
transform 1 0 74060 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_805
timestamp 1
transform 1 0 75164 0 1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_811
timestamp 1
transform 1 0 75716 0 1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_166_813
timestamp 1636968456
transform 1 0 75900 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_825
timestamp 1636968456
transform 1 0 77004 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_837
timestamp 1636968456
transform 1 0 78108 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_849
timestamp 1636968456
transform 1 0 79212 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_861
timestamp 1
transform 1 0 80316 0 1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_867
timestamp 1
transform 1 0 80868 0 1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_166_869
timestamp 1636968456
transform 1 0 81052 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_881
timestamp 1636968456
transform 1 0 82156 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_893
timestamp 1636968456
transform 1 0 83260 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_905
timestamp 1636968456
transform 1 0 84364 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_917
timestamp 1
transform 1 0 85468 0 1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_923
timestamp 1
transform 1 0 86020 0 1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_166_925
timestamp 1636968456
transform 1 0 86204 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_937
timestamp 1636968456
transform 1 0 87308 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_949
timestamp 1636968456
transform 1 0 88412 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_961
timestamp 1636968456
transform 1 0 89516 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_973
timestamp 1
transform 1 0 90620 0 1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_979
timestamp 1
transform 1 0 91172 0 1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_166_981
timestamp 1636968456
transform 1 0 91356 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_993
timestamp 1636968456
transform 1 0 92460 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_1005
timestamp 1636968456
transform 1 0 93564 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_1017
timestamp 1636968456
transform 1 0 94668 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_166_1029
timestamp 1
transform 1 0 95772 0 1 92480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_166_1035
timestamp 1
transform 1 0 96324 0 1 92480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_166_1037
timestamp 1636968456
transform 1 0 96508 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_1049
timestamp 1636968456
transform 1 0 97612 0 1 92480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_166_1061
timestamp 1636968456
transform 1 0 98716 0 1 92480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_166_1073
timestamp 1
transform 1 0 99820 0 1 92480
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_167_3
timestamp 1636968456
transform 1 0 1380 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_15
timestamp 1636968456
transform 1 0 2484 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_27
timestamp 1636968456
transform 1 0 3588 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_39
timestamp 1636968456
transform 1 0 4692 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_167_51
timestamp 1
transform 1 0 5796 0 -1 93568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_167_55
timestamp 1
transform 1 0 6164 0 -1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_167_57
timestamp 1636968456
transform 1 0 6348 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_69
timestamp 1636968456
transform 1 0 7452 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_81
timestamp 1636968456
transform 1 0 8556 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_93
timestamp 1636968456
transform 1 0 9660 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_167_105
timestamp 1
transform 1 0 10764 0 -1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_167_111
timestamp 1
transform 1 0 11316 0 -1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_167_113
timestamp 1636968456
transform 1 0 11500 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_125
timestamp 1636968456
transform 1 0 12604 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_137
timestamp 1636968456
transform 1 0 13708 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_149
timestamp 1636968456
transform 1 0 14812 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_167_161
timestamp 1
transform 1 0 15916 0 -1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_167_167
timestamp 1
transform 1 0 16468 0 -1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_167_169
timestamp 1636968456
transform 1 0 16652 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_181
timestamp 1636968456
transform 1 0 17756 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_193
timestamp 1636968456
transform 1 0 18860 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_205
timestamp 1636968456
transform 1 0 19964 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_167_217
timestamp 1
transform 1 0 21068 0 -1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_167_223
timestamp 1
transform 1 0 21620 0 -1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_167_225
timestamp 1636968456
transform 1 0 21804 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_237
timestamp 1636968456
transform 1 0 22908 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_249
timestamp 1636968456
transform 1 0 24012 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_261
timestamp 1636968456
transform 1 0 25116 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_167_273
timestamp 1
transform 1 0 26220 0 -1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_167_279
timestamp 1
transform 1 0 26772 0 -1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_167_281
timestamp 1636968456
transform 1 0 26956 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_293
timestamp 1636968456
transform 1 0 28060 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_305
timestamp 1636968456
transform 1 0 29164 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_317
timestamp 1636968456
transform 1 0 30268 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_167_329
timestamp 1
transform 1 0 31372 0 -1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_167_335
timestamp 1
transform 1 0 31924 0 -1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_167_337
timestamp 1636968456
transform 1 0 32108 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_349
timestamp 1636968456
transform 1 0 33212 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_361
timestamp 1636968456
transform 1 0 34316 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_373
timestamp 1636968456
transform 1 0 35420 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_167_385
timestamp 1
transform 1 0 36524 0 -1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_167_391
timestamp 1
transform 1 0 37076 0 -1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_167_393
timestamp 1636968456
transform 1 0 37260 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_405
timestamp 1636968456
transform 1 0 38364 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_417
timestamp 1636968456
transform 1 0 39468 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_429
timestamp 1636968456
transform 1 0 40572 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_167_441
timestamp 1
transform 1 0 41676 0 -1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_167_447
timestamp 1
transform 1 0 42228 0 -1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_167_449
timestamp 1636968456
transform 1 0 42412 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_461
timestamp 1636968456
transform 1 0 43516 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_473
timestamp 1636968456
transform 1 0 44620 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_485
timestamp 1636968456
transform 1 0 45724 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_167_497
timestamp 1
transform 1 0 46828 0 -1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_167_503
timestamp 1
transform 1 0 47380 0 -1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_167_505
timestamp 1636968456
transform 1 0 47564 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_517
timestamp 1636968456
transform 1 0 48668 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_529
timestamp 1636968456
transform 1 0 49772 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_541
timestamp 1636968456
transform 1 0 50876 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_167_553
timestamp 1
transform 1 0 51980 0 -1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_167_559
timestamp 1
transform 1 0 52532 0 -1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_167_561
timestamp 1636968456
transform 1 0 52716 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_573
timestamp 1636968456
transform 1 0 53820 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_585
timestamp 1636968456
transform 1 0 54924 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_597
timestamp 1636968456
transform 1 0 56028 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_167_609
timestamp 1
transform 1 0 57132 0 -1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_167_615
timestamp 1
transform 1 0 57684 0 -1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_167_617
timestamp 1636968456
transform 1 0 57868 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_629
timestamp 1636968456
transform 1 0 58972 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_641
timestamp 1636968456
transform 1 0 60076 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_653
timestamp 1636968456
transform 1 0 61180 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_167_665
timestamp 1
transform 1 0 62284 0 -1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_167_671
timestamp 1
transform 1 0 62836 0 -1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_167_673
timestamp 1636968456
transform 1 0 63020 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_685
timestamp 1636968456
transform 1 0 64124 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_697
timestamp 1636968456
transform 1 0 65228 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_709
timestamp 1636968456
transform 1 0 66332 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_167_721
timestamp 1
transform 1 0 67436 0 -1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_167_727
timestamp 1
transform 1 0 67988 0 -1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_167_729
timestamp 1636968456
transform 1 0 68172 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_741
timestamp 1636968456
transform 1 0 69276 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_753
timestamp 1636968456
transform 1 0 70380 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_765
timestamp 1636968456
transform 1 0 71484 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_167_777
timestamp 1
transform 1 0 72588 0 -1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_167_783
timestamp 1
transform 1 0 73140 0 -1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_167_785
timestamp 1636968456
transform 1 0 73324 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_797
timestamp 1636968456
transform 1 0 74428 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_809
timestamp 1636968456
transform 1 0 75532 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_821
timestamp 1636968456
transform 1 0 76636 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_167_833
timestamp 1
transform 1 0 77740 0 -1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_167_839
timestamp 1
transform 1 0 78292 0 -1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_167_841
timestamp 1636968456
transform 1 0 78476 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_853
timestamp 1636968456
transform 1 0 79580 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_865
timestamp 1636968456
transform 1 0 80684 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_877
timestamp 1636968456
transform 1 0 81788 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_167_889
timestamp 1
transform 1 0 82892 0 -1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_167_895
timestamp 1
transform 1 0 83444 0 -1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_167_897
timestamp 1636968456
transform 1 0 83628 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_909
timestamp 1636968456
transform 1 0 84732 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_921
timestamp 1636968456
transform 1 0 85836 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_933
timestamp 1636968456
transform 1 0 86940 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_167_945
timestamp 1
transform 1 0 88044 0 -1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_167_951
timestamp 1
transform 1 0 88596 0 -1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_167_953
timestamp 1636968456
transform 1 0 88780 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_965
timestamp 1636968456
transform 1 0 89884 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_977
timestamp 1636968456
transform 1 0 90988 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_989
timestamp 1636968456
transform 1 0 92092 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_167_1001
timestamp 1
transform 1 0 93196 0 -1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_167_1007
timestamp 1
transform 1 0 93748 0 -1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_167_1009
timestamp 1636968456
transform 1 0 93932 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_1021
timestamp 1636968456
transform 1 0 95036 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_1033
timestamp 1636968456
transform 1 0 96140 0 -1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_167_1045
timestamp 1636968456
transform 1 0 97244 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_167_1057
timestamp 1
transform 1 0 98348 0 -1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_167_1063
timestamp 1
transform 1 0 98900 0 -1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_167_1065
timestamp 1636968456
transform 1 0 99084 0 -1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_167_1077
timestamp 1
transform 1 0 100188 0 -1 93568
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_168_3
timestamp 1636968456
transform 1 0 1380 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_15
timestamp 1636968456
transform 1 0 2484 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_168_27
timestamp 1
transform 1 0 3588 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_29
timestamp 1636968456
transform 1 0 3772 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_41
timestamp 1636968456
transform 1 0 4876 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_53
timestamp 1636968456
transform 1 0 5980 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_65
timestamp 1636968456
transform 1 0 7084 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_77
timestamp 1
transform 1 0 8188 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_83
timestamp 1
transform 1 0 8740 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_85
timestamp 1636968456
transform 1 0 8924 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_97
timestamp 1636968456
transform 1 0 10028 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_109
timestamp 1636968456
transform 1 0 11132 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_121
timestamp 1636968456
transform 1 0 12236 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_133
timestamp 1
transform 1 0 13340 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_139
timestamp 1
transform 1 0 13892 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_141
timestamp 1636968456
transform 1 0 14076 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_153
timestamp 1636968456
transform 1 0 15180 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_165
timestamp 1636968456
transform 1 0 16284 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_177
timestamp 1636968456
transform 1 0 17388 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_189
timestamp 1
transform 1 0 18492 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_195
timestamp 1
transform 1 0 19044 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_197
timestamp 1636968456
transform 1 0 19228 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_209
timestamp 1636968456
transform 1 0 20332 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_221
timestamp 1636968456
transform 1 0 21436 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_233
timestamp 1636968456
transform 1 0 22540 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_245
timestamp 1
transform 1 0 23644 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_251
timestamp 1
transform 1 0 24196 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_253
timestamp 1636968456
transform 1 0 24380 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_265
timestamp 1636968456
transform 1 0 25484 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_277
timestamp 1636968456
transform 1 0 26588 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_289
timestamp 1636968456
transform 1 0 27692 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_301
timestamp 1
transform 1 0 28796 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_307
timestamp 1
transform 1 0 29348 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_309
timestamp 1636968456
transform 1 0 29532 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_321
timestamp 1636968456
transform 1 0 30636 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_333
timestamp 1636968456
transform 1 0 31740 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_345
timestamp 1636968456
transform 1 0 32844 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_357
timestamp 1
transform 1 0 33948 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_363
timestamp 1
transform 1 0 34500 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_365
timestamp 1636968456
transform 1 0 34684 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_377
timestamp 1636968456
transform 1 0 35788 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_389
timestamp 1636968456
transform 1 0 36892 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_401
timestamp 1636968456
transform 1 0 37996 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_413
timestamp 1
transform 1 0 39100 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_419
timestamp 1
transform 1 0 39652 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_421
timestamp 1636968456
transform 1 0 39836 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_433
timestamp 1636968456
transform 1 0 40940 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_445
timestamp 1636968456
transform 1 0 42044 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_457
timestamp 1636968456
transform 1 0 43148 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_469
timestamp 1
transform 1 0 44252 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_475
timestamp 1
transform 1 0 44804 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_477
timestamp 1636968456
transform 1 0 44988 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_489
timestamp 1636968456
transform 1 0 46092 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_501
timestamp 1636968456
transform 1 0 47196 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_513
timestamp 1636968456
transform 1 0 48300 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_525
timestamp 1
transform 1 0 49404 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_531
timestamp 1
transform 1 0 49956 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_533
timestamp 1636968456
transform 1 0 50140 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_545
timestamp 1636968456
transform 1 0 51244 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_557
timestamp 1636968456
transform 1 0 52348 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_569
timestamp 1636968456
transform 1 0 53452 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_581
timestamp 1
transform 1 0 54556 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_587
timestamp 1
transform 1 0 55108 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_589
timestamp 1636968456
transform 1 0 55292 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_601
timestamp 1636968456
transform 1 0 56396 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_613
timestamp 1636968456
transform 1 0 57500 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_625
timestamp 1636968456
transform 1 0 58604 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_637
timestamp 1
transform 1 0 59708 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_643
timestamp 1
transform 1 0 60260 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_645
timestamp 1636968456
transform 1 0 60444 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_657
timestamp 1636968456
transform 1 0 61548 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_669
timestamp 1636968456
transform 1 0 62652 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_681
timestamp 1636968456
transform 1 0 63756 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_693
timestamp 1
transform 1 0 64860 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_699
timestamp 1
transform 1 0 65412 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_701
timestamp 1636968456
transform 1 0 65596 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_713
timestamp 1636968456
transform 1 0 66700 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_725
timestamp 1636968456
transform 1 0 67804 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_737
timestamp 1636968456
transform 1 0 68908 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_749
timestamp 1
transform 1 0 70012 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_755
timestamp 1
transform 1 0 70564 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_757
timestamp 1636968456
transform 1 0 70748 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_769
timestamp 1636968456
transform 1 0 71852 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_781
timestamp 1636968456
transform 1 0 72956 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_793
timestamp 1636968456
transform 1 0 74060 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_805
timestamp 1
transform 1 0 75164 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_811
timestamp 1
transform 1 0 75716 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_813
timestamp 1636968456
transform 1 0 75900 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_825
timestamp 1636968456
transform 1 0 77004 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_837
timestamp 1636968456
transform 1 0 78108 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_849
timestamp 1636968456
transform 1 0 79212 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_861
timestamp 1
transform 1 0 80316 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_867
timestamp 1
transform 1 0 80868 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_869
timestamp 1636968456
transform 1 0 81052 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_881
timestamp 1636968456
transform 1 0 82156 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_893
timestamp 1636968456
transform 1 0 83260 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_905
timestamp 1636968456
transform 1 0 84364 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_917
timestamp 1
transform 1 0 85468 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_923
timestamp 1
transform 1 0 86020 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_925
timestamp 1636968456
transform 1 0 86204 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_937
timestamp 1636968456
transform 1 0 87308 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_949
timestamp 1636968456
transform 1 0 88412 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_961
timestamp 1636968456
transform 1 0 89516 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_973
timestamp 1
transform 1 0 90620 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_979
timestamp 1
transform 1 0 91172 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_981
timestamp 1636968456
transform 1 0 91356 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_993
timestamp 1636968456
transform 1 0 92460 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_1005
timestamp 1636968456
transform 1 0 93564 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_1017
timestamp 1636968456
transform 1 0 94668 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_168_1029
timestamp 1
transform 1 0 95772 0 1 93568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_168_1035
timestamp 1
transform 1 0 96324 0 1 93568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_168_1037
timestamp 1636968456
transform 1 0 96508 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_1049
timestamp 1636968456
transform 1 0 97612 0 1 93568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_168_1061
timestamp 1636968456
transform 1 0 98716 0 1 93568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_168_1073
timestamp 1
transform 1 0 99820 0 1 93568
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_169_3
timestamp 1636968456
transform 1 0 1380 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_15
timestamp 1636968456
transform 1 0 2484 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_27
timestamp 1636968456
transform 1 0 3588 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_39
timestamp 1636968456
transform 1 0 4692 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_169_51
timestamp 1
transform 1 0 5796 0 -1 94656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_169_55
timestamp 1
transform 1 0 6164 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_57
timestamp 1636968456
transform 1 0 6348 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_69
timestamp 1636968456
transform 1 0 7452 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_81
timestamp 1636968456
transform 1 0 8556 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_93
timestamp 1636968456
transform 1 0 9660 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_105
timestamp 1
transform 1 0 10764 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_111
timestamp 1
transform 1 0 11316 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_113
timestamp 1636968456
transform 1 0 11500 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_125
timestamp 1636968456
transform 1 0 12604 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_137
timestamp 1636968456
transform 1 0 13708 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_149
timestamp 1636968456
transform 1 0 14812 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_161
timestamp 1
transform 1 0 15916 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_167
timestamp 1
transform 1 0 16468 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_169
timestamp 1636968456
transform 1 0 16652 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_181
timestamp 1636968456
transform 1 0 17756 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_193
timestamp 1636968456
transform 1 0 18860 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_205
timestamp 1636968456
transform 1 0 19964 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_217
timestamp 1
transform 1 0 21068 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_223
timestamp 1
transform 1 0 21620 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_225
timestamp 1636968456
transform 1 0 21804 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_237
timestamp 1636968456
transform 1 0 22908 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_249
timestamp 1636968456
transform 1 0 24012 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_261
timestamp 1636968456
transform 1 0 25116 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_273
timestamp 1
transform 1 0 26220 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_279
timestamp 1
transform 1 0 26772 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_281
timestamp 1636968456
transform 1 0 26956 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_293
timestamp 1636968456
transform 1 0 28060 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_305
timestamp 1636968456
transform 1 0 29164 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_317
timestamp 1636968456
transform 1 0 30268 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_329
timestamp 1
transform 1 0 31372 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_335
timestamp 1
transform 1 0 31924 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_337
timestamp 1636968456
transform 1 0 32108 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_349
timestamp 1636968456
transform 1 0 33212 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_361
timestamp 1636968456
transform 1 0 34316 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_373
timestamp 1636968456
transform 1 0 35420 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_385
timestamp 1
transform 1 0 36524 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_391
timestamp 1
transform 1 0 37076 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_393
timestamp 1636968456
transform 1 0 37260 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_405
timestamp 1636968456
transform 1 0 38364 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_417
timestamp 1636968456
transform 1 0 39468 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_429
timestamp 1636968456
transform 1 0 40572 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_441
timestamp 1
transform 1 0 41676 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_447
timestamp 1
transform 1 0 42228 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_449
timestamp 1636968456
transform 1 0 42412 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_461
timestamp 1636968456
transform 1 0 43516 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_473
timestamp 1636968456
transform 1 0 44620 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_485
timestamp 1636968456
transform 1 0 45724 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_497
timestamp 1
transform 1 0 46828 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_503
timestamp 1
transform 1 0 47380 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_505
timestamp 1636968456
transform 1 0 47564 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_517
timestamp 1636968456
transform 1 0 48668 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_529
timestamp 1636968456
transform 1 0 49772 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_541
timestamp 1636968456
transform 1 0 50876 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_553
timestamp 1
transform 1 0 51980 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_559
timestamp 1
transform 1 0 52532 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_561
timestamp 1636968456
transform 1 0 52716 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_573
timestamp 1636968456
transform 1 0 53820 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_585
timestamp 1636968456
transform 1 0 54924 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_597
timestamp 1636968456
transform 1 0 56028 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_609
timestamp 1
transform 1 0 57132 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_615
timestamp 1
transform 1 0 57684 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_617
timestamp 1636968456
transform 1 0 57868 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_629
timestamp 1636968456
transform 1 0 58972 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_641
timestamp 1636968456
transform 1 0 60076 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_653
timestamp 1636968456
transform 1 0 61180 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_665
timestamp 1
transform 1 0 62284 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_671
timestamp 1
transform 1 0 62836 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_673
timestamp 1636968456
transform 1 0 63020 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_685
timestamp 1636968456
transform 1 0 64124 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_697
timestamp 1636968456
transform 1 0 65228 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_709
timestamp 1636968456
transform 1 0 66332 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_721
timestamp 1
transform 1 0 67436 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_727
timestamp 1
transform 1 0 67988 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_729
timestamp 1636968456
transform 1 0 68172 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_741
timestamp 1636968456
transform 1 0 69276 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_753
timestamp 1636968456
transform 1 0 70380 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_765
timestamp 1636968456
transform 1 0 71484 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_777
timestamp 1
transform 1 0 72588 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_783
timestamp 1
transform 1 0 73140 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_785
timestamp 1636968456
transform 1 0 73324 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_797
timestamp 1636968456
transform 1 0 74428 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_809
timestamp 1636968456
transform 1 0 75532 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_821
timestamp 1636968456
transform 1 0 76636 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_833
timestamp 1
transform 1 0 77740 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_839
timestamp 1
transform 1 0 78292 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_841
timestamp 1636968456
transform 1 0 78476 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_853
timestamp 1636968456
transform 1 0 79580 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_865
timestamp 1636968456
transform 1 0 80684 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_877
timestamp 1636968456
transform 1 0 81788 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_889
timestamp 1
transform 1 0 82892 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_895
timestamp 1
transform 1 0 83444 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_897
timestamp 1636968456
transform 1 0 83628 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_909
timestamp 1636968456
transform 1 0 84732 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_921
timestamp 1636968456
transform 1 0 85836 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_933
timestamp 1636968456
transform 1 0 86940 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_945
timestamp 1
transform 1 0 88044 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_951
timestamp 1
transform 1 0 88596 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_953
timestamp 1636968456
transform 1 0 88780 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_965
timestamp 1636968456
transform 1 0 89884 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_977
timestamp 1636968456
transform 1 0 90988 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_989
timestamp 1636968456
transform 1 0 92092 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_1001
timestamp 1
transform 1 0 93196 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_1007
timestamp 1
transform 1 0 93748 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_1009
timestamp 1636968456
transform 1 0 93932 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_1021
timestamp 1636968456
transform 1 0 95036 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_1033
timestamp 1636968456
transform 1 0 96140 0 -1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_169_1045
timestamp 1636968456
transform 1 0 97244 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_169_1057
timestamp 1
transform 1 0 98348 0 -1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_169_1063
timestamp 1
transform 1 0 98900 0 -1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_169_1065
timestamp 1636968456
transform 1 0 99084 0 -1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_169_1077
timestamp 1
transform 1 0 100188 0 -1 94656
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_170_3
timestamp 1636968456
transform 1 0 1380 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_15
timestamp 1636968456
transform 1 0 2484 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_170_27
timestamp 1
transform 1 0 3588 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_29
timestamp 1636968456
transform 1 0 3772 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_41
timestamp 1636968456
transform 1 0 4876 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_53
timestamp 1636968456
transform 1 0 5980 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_65
timestamp 1636968456
transform 1 0 7084 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_77
timestamp 1
transform 1 0 8188 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_83
timestamp 1
transform 1 0 8740 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_85
timestamp 1636968456
transform 1 0 8924 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_97
timestamp 1636968456
transform 1 0 10028 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_109
timestamp 1636968456
transform 1 0 11132 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_121
timestamp 1636968456
transform 1 0 12236 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_133
timestamp 1
transform 1 0 13340 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_139
timestamp 1
transform 1 0 13892 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_141
timestamp 1636968456
transform 1 0 14076 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_153
timestamp 1636968456
transform 1 0 15180 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_165
timestamp 1636968456
transform 1 0 16284 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_177
timestamp 1636968456
transform 1 0 17388 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_189
timestamp 1
transform 1 0 18492 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_195
timestamp 1
transform 1 0 19044 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_197
timestamp 1636968456
transform 1 0 19228 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_209
timestamp 1636968456
transform 1 0 20332 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_221
timestamp 1636968456
transform 1 0 21436 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_233
timestamp 1636968456
transform 1 0 22540 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_245
timestamp 1
transform 1 0 23644 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_251
timestamp 1
transform 1 0 24196 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_253
timestamp 1636968456
transform 1 0 24380 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_265
timestamp 1636968456
transform 1 0 25484 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_277
timestamp 1636968456
transform 1 0 26588 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_289
timestamp 1636968456
transform 1 0 27692 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_301
timestamp 1
transform 1 0 28796 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_307
timestamp 1
transform 1 0 29348 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_309
timestamp 1636968456
transform 1 0 29532 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_321
timestamp 1636968456
transform 1 0 30636 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_333
timestamp 1636968456
transform 1 0 31740 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_345
timestamp 1636968456
transform 1 0 32844 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_357
timestamp 1
transform 1 0 33948 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_363
timestamp 1
transform 1 0 34500 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_365
timestamp 1636968456
transform 1 0 34684 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_377
timestamp 1636968456
transform 1 0 35788 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_389
timestamp 1636968456
transform 1 0 36892 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_401
timestamp 1636968456
transform 1 0 37996 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_413
timestamp 1
transform 1 0 39100 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_419
timestamp 1
transform 1 0 39652 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_421
timestamp 1636968456
transform 1 0 39836 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_433
timestamp 1636968456
transform 1 0 40940 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_445
timestamp 1636968456
transform 1 0 42044 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_457
timestamp 1636968456
transform 1 0 43148 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_469
timestamp 1
transform 1 0 44252 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_475
timestamp 1
transform 1 0 44804 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_477
timestamp 1636968456
transform 1 0 44988 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_489
timestamp 1636968456
transform 1 0 46092 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_501
timestamp 1636968456
transform 1 0 47196 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_513
timestamp 1636968456
transform 1 0 48300 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_525
timestamp 1
transform 1 0 49404 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_531
timestamp 1
transform 1 0 49956 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_533
timestamp 1636968456
transform 1 0 50140 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_545
timestamp 1636968456
transform 1 0 51244 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_557
timestamp 1636968456
transform 1 0 52348 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_569
timestamp 1636968456
transform 1 0 53452 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_581
timestamp 1
transform 1 0 54556 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_587
timestamp 1
transform 1 0 55108 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_589
timestamp 1636968456
transform 1 0 55292 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_601
timestamp 1636968456
transform 1 0 56396 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_613
timestamp 1636968456
transform 1 0 57500 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_625
timestamp 1636968456
transform 1 0 58604 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_637
timestamp 1
transform 1 0 59708 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_643
timestamp 1
transform 1 0 60260 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_645
timestamp 1636968456
transform 1 0 60444 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_657
timestamp 1636968456
transform 1 0 61548 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_669
timestamp 1636968456
transform 1 0 62652 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_681
timestamp 1636968456
transform 1 0 63756 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_693
timestamp 1
transform 1 0 64860 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_699
timestamp 1
transform 1 0 65412 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_701
timestamp 1636968456
transform 1 0 65596 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_713
timestamp 1636968456
transform 1 0 66700 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_725
timestamp 1636968456
transform 1 0 67804 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_737
timestamp 1636968456
transform 1 0 68908 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_749
timestamp 1
transform 1 0 70012 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_755
timestamp 1
transform 1 0 70564 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_757
timestamp 1636968456
transform 1 0 70748 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_769
timestamp 1636968456
transform 1 0 71852 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_781
timestamp 1636968456
transform 1 0 72956 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_793
timestamp 1636968456
transform 1 0 74060 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_805
timestamp 1
transform 1 0 75164 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_811
timestamp 1
transform 1 0 75716 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_813
timestamp 1636968456
transform 1 0 75900 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_825
timestamp 1636968456
transform 1 0 77004 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_837
timestamp 1636968456
transform 1 0 78108 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_849
timestamp 1636968456
transform 1 0 79212 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_861
timestamp 1
transform 1 0 80316 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_867
timestamp 1
transform 1 0 80868 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_869
timestamp 1636968456
transform 1 0 81052 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_881
timestamp 1636968456
transform 1 0 82156 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_893
timestamp 1636968456
transform 1 0 83260 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_905
timestamp 1636968456
transform 1 0 84364 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_917
timestamp 1
transform 1 0 85468 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_923
timestamp 1
transform 1 0 86020 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_925
timestamp 1636968456
transform 1 0 86204 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_937
timestamp 1636968456
transform 1 0 87308 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_949
timestamp 1636968456
transform 1 0 88412 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_961
timestamp 1636968456
transform 1 0 89516 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_973
timestamp 1
transform 1 0 90620 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_979
timestamp 1
transform 1 0 91172 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_981
timestamp 1636968456
transform 1 0 91356 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_993
timestamp 1636968456
transform 1 0 92460 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_1005
timestamp 1636968456
transform 1 0 93564 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_1017
timestamp 1636968456
transform 1 0 94668 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_170_1029
timestamp 1
transform 1 0 95772 0 1 94656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_170_1035
timestamp 1
transform 1 0 96324 0 1 94656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_170_1037
timestamp 1636968456
transform 1 0 96508 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_1049
timestamp 1636968456
transform 1 0 97612 0 1 94656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_170_1061
timestamp 1636968456
transform 1 0 98716 0 1 94656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_170_1073
timestamp 1
transform 1 0 99820 0 1 94656
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_171_3
timestamp 1636968456
transform 1 0 1380 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_15
timestamp 1636968456
transform 1 0 2484 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_27
timestamp 1636968456
transform 1 0 3588 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_39
timestamp 1636968456
transform 1 0 4692 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_171_51
timestamp 1
transform 1 0 5796 0 -1 95744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_171_55
timestamp 1
transform 1 0 6164 0 -1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_171_57
timestamp 1636968456
transform 1 0 6348 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_69
timestamp 1636968456
transform 1 0 7452 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_81
timestamp 1636968456
transform 1 0 8556 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_93
timestamp 1636968456
transform 1 0 9660 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_171_105
timestamp 1
transform 1 0 10764 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_111
timestamp 1
transform 1 0 11316 0 -1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_171_113
timestamp 1636968456
transform 1 0 11500 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_125
timestamp 1636968456
transform 1 0 12604 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_137
timestamp 1636968456
transform 1 0 13708 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_149
timestamp 1636968456
transform 1 0 14812 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_171_161
timestamp 1
transform 1 0 15916 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_167
timestamp 1
transform 1 0 16468 0 -1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_171_169
timestamp 1636968456
transform 1 0 16652 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_181
timestamp 1636968456
transform 1 0 17756 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_193
timestamp 1636968456
transform 1 0 18860 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_205
timestamp 1636968456
transform 1 0 19964 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_171_217
timestamp 1
transform 1 0 21068 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_223
timestamp 1
transform 1 0 21620 0 -1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_171_225
timestamp 1636968456
transform 1 0 21804 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_237
timestamp 1636968456
transform 1 0 22908 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_249
timestamp 1636968456
transform 1 0 24012 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_261
timestamp 1636968456
transform 1 0 25116 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_171_273
timestamp 1
transform 1 0 26220 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_279
timestamp 1
transform 1 0 26772 0 -1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_171_281
timestamp 1636968456
transform 1 0 26956 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_293
timestamp 1636968456
transform 1 0 28060 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_305
timestamp 1636968456
transform 1 0 29164 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_317
timestamp 1636968456
transform 1 0 30268 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_171_329
timestamp 1
transform 1 0 31372 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_335
timestamp 1
transform 1 0 31924 0 -1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_171_337
timestamp 1636968456
transform 1 0 32108 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_349
timestamp 1636968456
transform 1 0 33212 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_361
timestamp 1636968456
transform 1 0 34316 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_373
timestamp 1636968456
transform 1 0 35420 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_171_385
timestamp 1
transform 1 0 36524 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_391
timestamp 1
transform 1 0 37076 0 -1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_171_393
timestamp 1636968456
transform 1 0 37260 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_405
timestamp 1636968456
transform 1 0 38364 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_417
timestamp 1636968456
transform 1 0 39468 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_429
timestamp 1636968456
transform 1 0 40572 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_171_441
timestamp 1
transform 1 0 41676 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_447
timestamp 1
transform 1 0 42228 0 -1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_171_449
timestamp 1636968456
transform 1 0 42412 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_461
timestamp 1636968456
transform 1 0 43516 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_473
timestamp 1636968456
transform 1 0 44620 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_485
timestamp 1636968456
transform 1 0 45724 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_171_497
timestamp 1
transform 1 0 46828 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_503
timestamp 1
transform 1 0 47380 0 -1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_171_505
timestamp 1636968456
transform 1 0 47564 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_517
timestamp 1636968456
transform 1 0 48668 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_529
timestamp 1636968456
transform 1 0 49772 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_541
timestamp 1636968456
transform 1 0 50876 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_171_553
timestamp 1
transform 1 0 51980 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_559
timestamp 1
transform 1 0 52532 0 -1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_171_561
timestamp 1636968456
transform 1 0 52716 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_573
timestamp 1636968456
transform 1 0 53820 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_585
timestamp 1636968456
transform 1 0 54924 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_597
timestamp 1636968456
transform 1 0 56028 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_171_609
timestamp 1
transform 1 0 57132 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_615
timestamp 1
transform 1 0 57684 0 -1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_171_617
timestamp 1636968456
transform 1 0 57868 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_629
timestamp 1636968456
transform 1 0 58972 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_641
timestamp 1636968456
transform 1 0 60076 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_653
timestamp 1636968456
transform 1 0 61180 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_171_665
timestamp 1
transform 1 0 62284 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_671
timestamp 1
transform 1 0 62836 0 -1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_171_673
timestamp 1636968456
transform 1 0 63020 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_685
timestamp 1636968456
transform 1 0 64124 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_697
timestamp 1636968456
transform 1 0 65228 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_709
timestamp 1636968456
transform 1 0 66332 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_171_721
timestamp 1
transform 1 0 67436 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_727
timestamp 1
transform 1 0 67988 0 -1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_171_729
timestamp 1636968456
transform 1 0 68172 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_741
timestamp 1636968456
transform 1 0 69276 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_753
timestamp 1636968456
transform 1 0 70380 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_765
timestamp 1636968456
transform 1 0 71484 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_171_777
timestamp 1
transform 1 0 72588 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_783
timestamp 1
transform 1 0 73140 0 -1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_171_785
timestamp 1636968456
transform 1 0 73324 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_797
timestamp 1636968456
transform 1 0 74428 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_809
timestamp 1636968456
transform 1 0 75532 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_821
timestamp 1636968456
transform 1 0 76636 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_171_833
timestamp 1
transform 1 0 77740 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_839
timestamp 1
transform 1 0 78292 0 -1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_171_841
timestamp 1636968456
transform 1 0 78476 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_853
timestamp 1636968456
transform 1 0 79580 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_865
timestamp 1636968456
transform 1 0 80684 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_877
timestamp 1636968456
transform 1 0 81788 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_171_889
timestamp 1
transform 1 0 82892 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_895
timestamp 1
transform 1 0 83444 0 -1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_171_897
timestamp 1636968456
transform 1 0 83628 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_909
timestamp 1636968456
transform 1 0 84732 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_921
timestamp 1636968456
transform 1 0 85836 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_933
timestamp 1636968456
transform 1 0 86940 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_171_945
timestamp 1
transform 1 0 88044 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_951
timestamp 1
transform 1 0 88596 0 -1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_171_953
timestamp 1636968456
transform 1 0 88780 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_965
timestamp 1636968456
transform 1 0 89884 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_977
timestamp 1636968456
transform 1 0 90988 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_989
timestamp 1636968456
transform 1 0 92092 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_171_1001
timestamp 1
transform 1 0 93196 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_1007
timestamp 1
transform 1 0 93748 0 -1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_171_1009
timestamp 1636968456
transform 1 0 93932 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_1021
timestamp 1636968456
transform 1 0 95036 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_1033
timestamp 1636968456
transform 1 0 96140 0 -1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_171_1045
timestamp 1636968456
transform 1 0 97244 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_171_1057
timestamp 1
transform 1 0 98348 0 -1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_171_1063
timestamp 1
transform 1 0 98900 0 -1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_171_1065
timestamp 1636968456
transform 1 0 99084 0 -1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_171_1077
timestamp 1
transform 1 0 100188 0 -1 95744
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_172_3
timestamp 1636968456
transform 1 0 1380 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_15
timestamp 1636968456
transform 1 0 2484 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_172_27
timestamp 1
transform 1 0 3588 0 1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_172_29
timestamp 1636968456
transform 1 0 3772 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_41
timestamp 1636968456
transform 1 0 4876 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_53
timestamp 1636968456
transform 1 0 5980 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_65
timestamp 1636968456
transform 1 0 7084 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_172_77
timestamp 1
transform 1 0 8188 0 1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_172_83
timestamp 1
transform 1 0 8740 0 1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_172_85
timestamp 1636968456
transform 1 0 8924 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_97
timestamp 1636968456
transform 1 0 10028 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_109
timestamp 1636968456
transform 1 0 11132 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_121
timestamp 1636968456
transform 1 0 12236 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_172_133
timestamp 1
transform 1 0 13340 0 1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_172_139
timestamp 1
transform 1 0 13892 0 1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_172_141
timestamp 1636968456
transform 1 0 14076 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_153
timestamp 1636968456
transform 1 0 15180 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_165
timestamp 1636968456
transform 1 0 16284 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_177
timestamp 1636968456
transform 1 0 17388 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_172_189
timestamp 1
transform 1 0 18492 0 1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_172_195
timestamp 1
transform 1 0 19044 0 1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_172_197
timestamp 1636968456
transform 1 0 19228 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_209
timestamp 1636968456
transform 1 0 20332 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_221
timestamp 1636968456
transform 1 0 21436 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_233
timestamp 1636968456
transform 1 0 22540 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_172_245
timestamp 1
transform 1 0 23644 0 1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_172_251
timestamp 1
transform 1 0 24196 0 1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_172_253
timestamp 1636968456
transform 1 0 24380 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_265
timestamp 1636968456
transform 1 0 25484 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_277
timestamp 1636968456
transform 1 0 26588 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_289
timestamp 1636968456
transform 1 0 27692 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_172_301
timestamp 1
transform 1 0 28796 0 1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_172_307
timestamp 1
transform 1 0 29348 0 1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_172_309
timestamp 1636968456
transform 1 0 29532 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_321
timestamp 1636968456
transform 1 0 30636 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_333
timestamp 1636968456
transform 1 0 31740 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_345
timestamp 1636968456
transform 1 0 32844 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_172_357
timestamp 1
transform 1 0 33948 0 1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_172_363
timestamp 1
transform 1 0 34500 0 1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_172_365
timestamp 1636968456
transform 1 0 34684 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_377
timestamp 1636968456
transform 1 0 35788 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_389
timestamp 1636968456
transform 1 0 36892 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_401
timestamp 1636968456
transform 1 0 37996 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_172_413
timestamp 1
transform 1 0 39100 0 1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_172_419
timestamp 1
transform 1 0 39652 0 1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_172_421
timestamp 1636968456
transform 1 0 39836 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_433
timestamp 1636968456
transform 1 0 40940 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_445
timestamp 1636968456
transform 1 0 42044 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_457
timestamp 1636968456
transform 1 0 43148 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_172_469
timestamp 1
transform 1 0 44252 0 1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_172_475
timestamp 1
transform 1 0 44804 0 1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_172_477
timestamp 1636968456
transform 1 0 44988 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_489
timestamp 1636968456
transform 1 0 46092 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_501
timestamp 1636968456
transform 1 0 47196 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_513
timestamp 1636968456
transform 1 0 48300 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_172_525
timestamp 1
transform 1 0 49404 0 1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_172_531
timestamp 1
transform 1 0 49956 0 1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_172_533
timestamp 1636968456
transform 1 0 50140 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_545
timestamp 1636968456
transform 1 0 51244 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_557
timestamp 1636968456
transform 1 0 52348 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_569
timestamp 1636968456
transform 1 0 53452 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_172_581
timestamp 1
transform 1 0 54556 0 1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_172_587
timestamp 1
transform 1 0 55108 0 1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_172_589
timestamp 1636968456
transform 1 0 55292 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_601
timestamp 1636968456
transform 1 0 56396 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_613
timestamp 1636968456
transform 1 0 57500 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_625
timestamp 1636968456
transform 1 0 58604 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_172_637
timestamp 1
transform 1 0 59708 0 1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_172_643
timestamp 1
transform 1 0 60260 0 1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_172_645
timestamp 1636968456
transform 1 0 60444 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_657
timestamp 1636968456
transform 1 0 61548 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_669
timestamp 1636968456
transform 1 0 62652 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_681
timestamp 1636968456
transform 1 0 63756 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_172_693
timestamp 1
transform 1 0 64860 0 1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_172_699
timestamp 1
transform 1 0 65412 0 1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_172_701
timestamp 1636968456
transform 1 0 65596 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_713
timestamp 1636968456
transform 1 0 66700 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_725
timestamp 1636968456
transform 1 0 67804 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_737
timestamp 1636968456
transform 1 0 68908 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_172_749
timestamp 1
transform 1 0 70012 0 1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_172_755
timestamp 1
transform 1 0 70564 0 1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_172_757
timestamp 1636968456
transform 1 0 70748 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_769
timestamp 1636968456
transform 1 0 71852 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_781
timestamp 1636968456
transform 1 0 72956 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_793
timestamp 1636968456
transform 1 0 74060 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_172_805
timestamp 1
transform 1 0 75164 0 1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_172_811
timestamp 1
transform 1 0 75716 0 1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_172_813
timestamp 1636968456
transform 1 0 75900 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_825
timestamp 1636968456
transform 1 0 77004 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_837
timestamp 1636968456
transform 1 0 78108 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_849
timestamp 1636968456
transform 1 0 79212 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_172_861
timestamp 1
transform 1 0 80316 0 1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_172_867
timestamp 1
transform 1 0 80868 0 1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_172_869
timestamp 1636968456
transform 1 0 81052 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_881
timestamp 1636968456
transform 1 0 82156 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_893
timestamp 1636968456
transform 1 0 83260 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_905
timestamp 1636968456
transform 1 0 84364 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_172_917
timestamp 1
transform 1 0 85468 0 1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_172_923
timestamp 1
transform 1 0 86020 0 1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_172_925
timestamp 1636968456
transform 1 0 86204 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_937
timestamp 1636968456
transform 1 0 87308 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_949
timestamp 1636968456
transform 1 0 88412 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_961
timestamp 1636968456
transform 1 0 89516 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_172_973
timestamp 1
transform 1 0 90620 0 1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_172_979
timestamp 1
transform 1 0 91172 0 1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_172_981
timestamp 1636968456
transform 1 0 91356 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_993
timestamp 1636968456
transform 1 0 92460 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_1005
timestamp 1636968456
transform 1 0 93564 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_1017
timestamp 1636968456
transform 1 0 94668 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_172_1029
timestamp 1
transform 1 0 95772 0 1 95744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_172_1035
timestamp 1
transform 1 0 96324 0 1 95744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_172_1037
timestamp 1636968456
transform 1 0 96508 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_1049
timestamp 1636968456
transform 1 0 97612 0 1 95744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_172_1061
timestamp 1636968456
transform 1 0 98716 0 1 95744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_172_1073
timestamp 1
transform 1 0 99820 0 1 95744
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_173_3
timestamp 1636968456
transform 1 0 1380 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_15
timestamp 1636968456
transform 1 0 2484 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_27
timestamp 1636968456
transform 1 0 3588 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_39
timestamp 1636968456
transform 1 0 4692 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_173_51
timestamp 1
transform 1 0 5796 0 -1 96832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_173_55
timestamp 1
transform 1 0 6164 0 -1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_173_57
timestamp 1636968456
transform 1 0 6348 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_69
timestamp 1636968456
transform 1 0 7452 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_81
timestamp 1636968456
transform 1 0 8556 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_93
timestamp 1636968456
transform 1 0 9660 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_173_105
timestamp 1
transform 1 0 10764 0 -1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_173_111
timestamp 1
transform 1 0 11316 0 -1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_173_113
timestamp 1636968456
transform 1 0 11500 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_125
timestamp 1636968456
transform 1 0 12604 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_137
timestamp 1636968456
transform 1 0 13708 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_149
timestamp 1636968456
transform 1 0 14812 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_173_161
timestamp 1
transform 1 0 15916 0 -1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_173_167
timestamp 1
transform 1 0 16468 0 -1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_173_169
timestamp 1636968456
transform 1 0 16652 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_181
timestamp 1636968456
transform 1 0 17756 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_193
timestamp 1636968456
transform 1 0 18860 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_205
timestamp 1636968456
transform 1 0 19964 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_173_217
timestamp 1
transform 1 0 21068 0 -1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_173_223
timestamp 1
transform 1 0 21620 0 -1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_173_225
timestamp 1636968456
transform 1 0 21804 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_237
timestamp 1636968456
transform 1 0 22908 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_249
timestamp 1636968456
transform 1 0 24012 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_261
timestamp 1636968456
transform 1 0 25116 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_173_273
timestamp 1
transform 1 0 26220 0 -1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_173_279
timestamp 1
transform 1 0 26772 0 -1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_173_281
timestamp 1636968456
transform 1 0 26956 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_293
timestamp 1636968456
transform 1 0 28060 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_305
timestamp 1636968456
transform 1 0 29164 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_317
timestamp 1636968456
transform 1 0 30268 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_173_329
timestamp 1
transform 1 0 31372 0 -1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_173_335
timestamp 1
transform 1 0 31924 0 -1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_173_337
timestamp 1636968456
transform 1 0 32108 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_349
timestamp 1636968456
transform 1 0 33212 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_361
timestamp 1636968456
transform 1 0 34316 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_373
timestamp 1636968456
transform 1 0 35420 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_173_385
timestamp 1
transform 1 0 36524 0 -1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_173_391
timestamp 1
transform 1 0 37076 0 -1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_173_393
timestamp 1636968456
transform 1 0 37260 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_405
timestamp 1636968456
transform 1 0 38364 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_417
timestamp 1636968456
transform 1 0 39468 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_429
timestamp 1636968456
transform 1 0 40572 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_173_441
timestamp 1
transform 1 0 41676 0 -1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_173_447
timestamp 1
transform 1 0 42228 0 -1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_173_449
timestamp 1636968456
transform 1 0 42412 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_461
timestamp 1636968456
transform 1 0 43516 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_473
timestamp 1636968456
transform 1 0 44620 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_485
timestamp 1636968456
transform 1 0 45724 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_173_497
timestamp 1
transform 1 0 46828 0 -1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_173_503
timestamp 1
transform 1 0 47380 0 -1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_173_505
timestamp 1636968456
transform 1 0 47564 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_517
timestamp 1636968456
transform 1 0 48668 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_529
timestamp 1636968456
transform 1 0 49772 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_541
timestamp 1636968456
transform 1 0 50876 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_173_553
timestamp 1
transform 1 0 51980 0 -1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_173_559
timestamp 1
transform 1 0 52532 0 -1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_173_561
timestamp 1636968456
transform 1 0 52716 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_573
timestamp 1636968456
transform 1 0 53820 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_585
timestamp 1636968456
transform 1 0 54924 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_597
timestamp 1636968456
transform 1 0 56028 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_173_609
timestamp 1
transform 1 0 57132 0 -1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_173_615
timestamp 1
transform 1 0 57684 0 -1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_173_617
timestamp 1636968456
transform 1 0 57868 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_629
timestamp 1636968456
transform 1 0 58972 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_641
timestamp 1636968456
transform 1 0 60076 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_653
timestamp 1636968456
transform 1 0 61180 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_173_665
timestamp 1
transform 1 0 62284 0 -1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_173_671
timestamp 1
transform 1 0 62836 0 -1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_173_673
timestamp 1636968456
transform 1 0 63020 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_685
timestamp 1636968456
transform 1 0 64124 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_697
timestamp 1636968456
transform 1 0 65228 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_709
timestamp 1636968456
transform 1 0 66332 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_173_721
timestamp 1
transform 1 0 67436 0 -1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_173_727
timestamp 1
transform 1 0 67988 0 -1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_173_729
timestamp 1636968456
transform 1 0 68172 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_741
timestamp 1636968456
transform 1 0 69276 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_753
timestamp 1636968456
transform 1 0 70380 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_765
timestamp 1636968456
transform 1 0 71484 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_173_777
timestamp 1
transform 1 0 72588 0 -1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_173_783
timestamp 1
transform 1 0 73140 0 -1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_173_785
timestamp 1636968456
transform 1 0 73324 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_797
timestamp 1636968456
transform 1 0 74428 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_809
timestamp 1636968456
transform 1 0 75532 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_821
timestamp 1636968456
transform 1 0 76636 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_173_833
timestamp 1
transform 1 0 77740 0 -1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_173_839
timestamp 1
transform 1 0 78292 0 -1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_173_841
timestamp 1636968456
transform 1 0 78476 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_853
timestamp 1636968456
transform 1 0 79580 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_865
timestamp 1636968456
transform 1 0 80684 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_877
timestamp 1636968456
transform 1 0 81788 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_173_889
timestamp 1
transform 1 0 82892 0 -1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_173_895
timestamp 1
transform 1 0 83444 0 -1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_173_897
timestamp 1636968456
transform 1 0 83628 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_909
timestamp 1636968456
transform 1 0 84732 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_921
timestamp 1636968456
transform 1 0 85836 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_933
timestamp 1636968456
transform 1 0 86940 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_173_945
timestamp 1
transform 1 0 88044 0 -1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_173_951
timestamp 1
transform 1 0 88596 0 -1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_173_953
timestamp 1636968456
transform 1 0 88780 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_965
timestamp 1636968456
transform 1 0 89884 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_977
timestamp 1636968456
transform 1 0 90988 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_989
timestamp 1636968456
transform 1 0 92092 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_173_1001
timestamp 1
transform 1 0 93196 0 -1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_173_1007
timestamp 1
transform 1 0 93748 0 -1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_173_1009
timestamp 1636968456
transform 1 0 93932 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_1021
timestamp 1636968456
transform 1 0 95036 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_1033
timestamp 1636968456
transform 1 0 96140 0 -1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_173_1045
timestamp 1636968456
transform 1 0 97244 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_173_1057
timestamp 1
transform 1 0 98348 0 -1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_173_1063
timestamp 1
transform 1 0 98900 0 -1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_173_1065
timestamp 1636968456
transform 1 0 99084 0 -1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_173_1077
timestamp 1
transform 1 0 100188 0 -1 96832
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_174_3
timestamp 1636968456
transform 1 0 1380 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_15
timestamp 1636968456
transform 1 0 2484 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_174_27
timestamp 1
transform 1 0 3588 0 1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_174_29
timestamp 1636968456
transform 1 0 3772 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_41
timestamp 1636968456
transform 1 0 4876 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_53
timestamp 1636968456
transform 1 0 5980 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_65
timestamp 1636968456
transform 1 0 7084 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_174_77
timestamp 1
transform 1 0 8188 0 1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_174_83
timestamp 1
transform 1 0 8740 0 1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_174_85
timestamp 1636968456
transform 1 0 8924 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_97
timestamp 1636968456
transform 1 0 10028 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_109
timestamp 1636968456
transform 1 0 11132 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_121
timestamp 1636968456
transform 1 0 12236 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_174_133
timestamp 1
transform 1 0 13340 0 1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_174_139
timestamp 1
transform 1 0 13892 0 1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_174_141
timestamp 1636968456
transform 1 0 14076 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_153
timestamp 1636968456
transform 1 0 15180 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_165
timestamp 1636968456
transform 1 0 16284 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_177
timestamp 1636968456
transform 1 0 17388 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_174_189
timestamp 1
transform 1 0 18492 0 1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_174_195
timestamp 1
transform 1 0 19044 0 1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_174_197
timestamp 1636968456
transform 1 0 19228 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_209
timestamp 1636968456
transform 1 0 20332 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_221
timestamp 1636968456
transform 1 0 21436 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_233
timestamp 1636968456
transform 1 0 22540 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_174_245
timestamp 1
transform 1 0 23644 0 1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_174_251
timestamp 1
transform 1 0 24196 0 1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_174_253
timestamp 1636968456
transform 1 0 24380 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_265
timestamp 1636968456
transform 1 0 25484 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_277
timestamp 1636968456
transform 1 0 26588 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_289
timestamp 1636968456
transform 1 0 27692 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_174_301
timestamp 1
transform 1 0 28796 0 1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_174_307
timestamp 1
transform 1 0 29348 0 1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_174_309
timestamp 1636968456
transform 1 0 29532 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_321
timestamp 1636968456
transform 1 0 30636 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_333
timestamp 1636968456
transform 1 0 31740 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_345
timestamp 1636968456
transform 1 0 32844 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_174_357
timestamp 1
transform 1 0 33948 0 1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_174_363
timestamp 1
transform 1 0 34500 0 1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_174_365
timestamp 1636968456
transform 1 0 34684 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_377
timestamp 1636968456
transform 1 0 35788 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_389
timestamp 1636968456
transform 1 0 36892 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_401
timestamp 1636968456
transform 1 0 37996 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_174_413
timestamp 1
transform 1 0 39100 0 1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_174_419
timestamp 1
transform 1 0 39652 0 1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_174_421
timestamp 1636968456
transform 1 0 39836 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_433
timestamp 1636968456
transform 1 0 40940 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_445
timestamp 1636968456
transform 1 0 42044 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_457
timestamp 1636968456
transform 1 0 43148 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_174_469
timestamp 1
transform 1 0 44252 0 1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_174_475
timestamp 1
transform 1 0 44804 0 1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_174_477
timestamp 1636968456
transform 1 0 44988 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_489
timestamp 1636968456
transform 1 0 46092 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_501
timestamp 1636968456
transform 1 0 47196 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_513
timestamp 1636968456
transform 1 0 48300 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_174_525
timestamp 1
transform 1 0 49404 0 1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_174_531
timestamp 1
transform 1 0 49956 0 1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_174_533
timestamp 1636968456
transform 1 0 50140 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_545
timestamp 1636968456
transform 1 0 51244 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_557
timestamp 1636968456
transform 1 0 52348 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_569
timestamp 1636968456
transform 1 0 53452 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_174_581
timestamp 1
transform 1 0 54556 0 1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_174_587
timestamp 1
transform 1 0 55108 0 1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_174_589
timestamp 1636968456
transform 1 0 55292 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_601
timestamp 1636968456
transform 1 0 56396 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_613
timestamp 1636968456
transform 1 0 57500 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_625
timestamp 1636968456
transform 1 0 58604 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_174_637
timestamp 1
transform 1 0 59708 0 1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_174_643
timestamp 1
transform 1 0 60260 0 1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_174_645
timestamp 1636968456
transform 1 0 60444 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_657
timestamp 1636968456
transform 1 0 61548 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_669
timestamp 1636968456
transform 1 0 62652 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_681
timestamp 1636968456
transform 1 0 63756 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_174_693
timestamp 1
transform 1 0 64860 0 1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_174_699
timestamp 1
transform 1 0 65412 0 1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_174_701
timestamp 1636968456
transform 1 0 65596 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_713
timestamp 1636968456
transform 1 0 66700 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_725
timestamp 1636968456
transform 1 0 67804 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_737
timestamp 1636968456
transform 1 0 68908 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_174_749
timestamp 1
transform 1 0 70012 0 1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_174_755
timestamp 1
transform 1 0 70564 0 1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_174_757
timestamp 1636968456
transform 1 0 70748 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_769
timestamp 1636968456
transform 1 0 71852 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_781
timestamp 1636968456
transform 1 0 72956 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_793
timestamp 1636968456
transform 1 0 74060 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_174_805
timestamp 1
transform 1 0 75164 0 1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_174_811
timestamp 1
transform 1 0 75716 0 1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_174_813
timestamp 1636968456
transform 1 0 75900 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_825
timestamp 1636968456
transform 1 0 77004 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_837
timestamp 1636968456
transform 1 0 78108 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_849
timestamp 1636968456
transform 1 0 79212 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_174_861
timestamp 1
transform 1 0 80316 0 1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_174_867
timestamp 1
transform 1 0 80868 0 1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_174_869
timestamp 1636968456
transform 1 0 81052 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_881
timestamp 1636968456
transform 1 0 82156 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_893
timestamp 1636968456
transform 1 0 83260 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_905
timestamp 1636968456
transform 1 0 84364 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_174_917
timestamp 1
transform 1 0 85468 0 1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_174_923
timestamp 1
transform 1 0 86020 0 1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_174_925
timestamp 1636968456
transform 1 0 86204 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_937
timestamp 1636968456
transform 1 0 87308 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_949
timestamp 1636968456
transform 1 0 88412 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_961
timestamp 1636968456
transform 1 0 89516 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_174_973
timestamp 1
transform 1 0 90620 0 1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_174_979
timestamp 1
transform 1 0 91172 0 1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_174_981
timestamp 1636968456
transform 1 0 91356 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_993
timestamp 1636968456
transform 1 0 92460 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_1005
timestamp 1636968456
transform 1 0 93564 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_1017
timestamp 1636968456
transform 1 0 94668 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_174_1029
timestamp 1
transform 1 0 95772 0 1 96832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_174_1035
timestamp 1
transform 1 0 96324 0 1 96832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_174_1037
timestamp 1636968456
transform 1 0 96508 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_1049
timestamp 1636968456
transform 1 0 97612 0 1 96832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_174_1061
timestamp 1636968456
transform 1 0 98716 0 1 96832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_174_1073
timestamp 1
transform 1 0 99820 0 1 96832
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_175_3
timestamp 1636968456
transform 1 0 1380 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_15
timestamp 1636968456
transform 1 0 2484 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_27
timestamp 1636968456
transform 1 0 3588 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_39
timestamp 1636968456
transform 1 0 4692 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_175_51
timestamp 1
transform 1 0 5796 0 -1 97920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_175_55
timestamp 1
transform 1 0 6164 0 -1 97920
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_175_57
timestamp 1636968456
transform 1 0 6348 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_69
timestamp 1636968456
transform 1 0 7452 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_81
timestamp 1636968456
transform 1 0 8556 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_93
timestamp 1636968456
transform 1 0 9660 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_175_105
timestamp 1
transform 1 0 10764 0 -1 97920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_175_111
timestamp 1
transform 1 0 11316 0 -1 97920
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_175_113
timestamp 1636968456
transform 1 0 11500 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_125
timestamp 1636968456
transform 1 0 12604 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_137
timestamp 1636968456
transform 1 0 13708 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_149
timestamp 1636968456
transform 1 0 14812 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_175_161
timestamp 1
transform 1 0 15916 0 -1 97920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_175_167
timestamp 1
transform 1 0 16468 0 -1 97920
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_175_169
timestamp 1636968456
transform 1 0 16652 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_181
timestamp 1636968456
transform 1 0 17756 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_193
timestamp 1636968456
transform 1 0 18860 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_205
timestamp 1636968456
transform 1 0 19964 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_175_217
timestamp 1
transform 1 0 21068 0 -1 97920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_175_223
timestamp 1
transform 1 0 21620 0 -1 97920
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_175_225
timestamp 1636968456
transform 1 0 21804 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_237
timestamp 1636968456
transform 1 0 22908 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_249
timestamp 1636968456
transform 1 0 24012 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_261
timestamp 1636968456
transform 1 0 25116 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_175_273
timestamp 1
transform 1 0 26220 0 -1 97920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_175_279
timestamp 1
transform 1 0 26772 0 -1 97920
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_175_281
timestamp 1636968456
transform 1 0 26956 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_293
timestamp 1636968456
transform 1 0 28060 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_305
timestamp 1636968456
transform 1 0 29164 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_317
timestamp 1636968456
transform 1 0 30268 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_175_329
timestamp 1
transform 1 0 31372 0 -1 97920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_175_335
timestamp 1
transform 1 0 31924 0 -1 97920
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_175_337
timestamp 1636968456
transform 1 0 32108 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_349
timestamp 1636968456
transform 1 0 33212 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_361
timestamp 1636968456
transform 1 0 34316 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_373
timestamp 1636968456
transform 1 0 35420 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_175_385
timestamp 1
transform 1 0 36524 0 -1 97920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_175_391
timestamp 1
transform 1 0 37076 0 -1 97920
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_175_393
timestamp 1636968456
transform 1 0 37260 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_405
timestamp 1636968456
transform 1 0 38364 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_417
timestamp 1636968456
transform 1 0 39468 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_429
timestamp 1636968456
transform 1 0 40572 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_175_441
timestamp 1
transform 1 0 41676 0 -1 97920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_175_447
timestamp 1
transform 1 0 42228 0 -1 97920
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_175_449
timestamp 1636968456
transform 1 0 42412 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_461
timestamp 1636968456
transform 1 0 43516 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_473
timestamp 1636968456
transform 1 0 44620 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_485
timestamp 1636968456
transform 1 0 45724 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_175_497
timestamp 1
transform 1 0 46828 0 -1 97920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_175_503
timestamp 1
transform 1 0 47380 0 -1 97920
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_175_505
timestamp 1636968456
transform 1 0 47564 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_517
timestamp 1636968456
transform 1 0 48668 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_529
timestamp 1636968456
transform 1 0 49772 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_541
timestamp 1636968456
transform 1 0 50876 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_175_553
timestamp 1
transform 1 0 51980 0 -1 97920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_175_559
timestamp 1
transform 1 0 52532 0 -1 97920
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_175_561
timestamp 1636968456
transform 1 0 52716 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_573
timestamp 1636968456
transform 1 0 53820 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_585
timestamp 1636968456
transform 1 0 54924 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_597
timestamp 1636968456
transform 1 0 56028 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_175_609
timestamp 1
transform 1 0 57132 0 -1 97920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_175_615
timestamp 1
transform 1 0 57684 0 -1 97920
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_175_617
timestamp 1636968456
transform 1 0 57868 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_629
timestamp 1636968456
transform 1 0 58972 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_641
timestamp 1636968456
transform 1 0 60076 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_653
timestamp 1636968456
transform 1 0 61180 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_175_665
timestamp 1
transform 1 0 62284 0 -1 97920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_175_671
timestamp 1
transform 1 0 62836 0 -1 97920
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_175_673
timestamp 1636968456
transform 1 0 63020 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_685
timestamp 1636968456
transform 1 0 64124 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_697
timestamp 1636968456
transform 1 0 65228 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_709
timestamp 1636968456
transform 1 0 66332 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_175_721
timestamp 1
transform 1 0 67436 0 -1 97920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_175_727
timestamp 1
transform 1 0 67988 0 -1 97920
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_175_729
timestamp 1636968456
transform 1 0 68172 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_741
timestamp 1636968456
transform 1 0 69276 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_753
timestamp 1636968456
transform 1 0 70380 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_765
timestamp 1636968456
transform 1 0 71484 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_175_777
timestamp 1
transform 1 0 72588 0 -1 97920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_175_783
timestamp 1
transform 1 0 73140 0 -1 97920
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_175_785
timestamp 1636968456
transform 1 0 73324 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_797
timestamp 1636968456
transform 1 0 74428 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_809
timestamp 1636968456
transform 1 0 75532 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_821
timestamp 1636968456
transform 1 0 76636 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_175_833
timestamp 1
transform 1 0 77740 0 -1 97920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_175_839
timestamp 1
transform 1 0 78292 0 -1 97920
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_175_841
timestamp 1636968456
transform 1 0 78476 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_853
timestamp 1636968456
transform 1 0 79580 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_865
timestamp 1636968456
transform 1 0 80684 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_877
timestamp 1636968456
transform 1 0 81788 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_175_889
timestamp 1
transform 1 0 82892 0 -1 97920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_175_895
timestamp 1
transform 1 0 83444 0 -1 97920
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_175_897
timestamp 1636968456
transform 1 0 83628 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_909
timestamp 1636968456
transform 1 0 84732 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_921
timestamp 1636968456
transform 1 0 85836 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_933
timestamp 1636968456
transform 1 0 86940 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_175_945
timestamp 1
transform 1 0 88044 0 -1 97920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_175_951
timestamp 1
transform 1 0 88596 0 -1 97920
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_175_953
timestamp 1636968456
transform 1 0 88780 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_965
timestamp 1636968456
transform 1 0 89884 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_977
timestamp 1636968456
transform 1 0 90988 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_989
timestamp 1636968456
transform 1 0 92092 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_175_1001
timestamp 1
transform 1 0 93196 0 -1 97920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_175_1007
timestamp 1
transform 1 0 93748 0 -1 97920
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_175_1009
timestamp 1636968456
transform 1 0 93932 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_1021
timestamp 1636968456
transform 1 0 95036 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_1033
timestamp 1636968456
transform 1 0 96140 0 -1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_175_1045
timestamp 1636968456
transform 1 0 97244 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_175_1057
timestamp 1
transform 1 0 98348 0 -1 97920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_175_1063
timestamp 1
transform 1 0 98900 0 -1 97920
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_175_1065
timestamp 1636968456
transform 1 0 99084 0 -1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_175_1077
timestamp 1
transform 1 0 100188 0 -1 97920
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_176_3
timestamp 1636968456
transform 1 0 1380 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_15
timestamp 1636968456
transform 1 0 2484 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_176_27
timestamp 1
transform 1 0 3588 0 1 97920
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_176_29
timestamp 1636968456
transform 1 0 3772 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_41
timestamp 1636968456
transform 1 0 4876 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_53
timestamp 1636968456
transform 1 0 5980 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_65
timestamp 1636968456
transform 1 0 7084 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_176_77
timestamp 1
transform 1 0 8188 0 1 97920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_176_83
timestamp 1
transform 1 0 8740 0 1 97920
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_176_85
timestamp 1636968456
transform 1 0 8924 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_97
timestamp 1636968456
transform 1 0 10028 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_109
timestamp 1636968456
transform 1 0 11132 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_121
timestamp 1636968456
transform 1 0 12236 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_176_133
timestamp 1
transform 1 0 13340 0 1 97920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_176_139
timestamp 1
transform 1 0 13892 0 1 97920
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_176_141
timestamp 1636968456
transform 1 0 14076 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_153
timestamp 1636968456
transform 1 0 15180 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_165
timestamp 1636968456
transform 1 0 16284 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_177
timestamp 1636968456
transform 1 0 17388 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_176_189
timestamp 1
transform 1 0 18492 0 1 97920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_176_195
timestamp 1
transform 1 0 19044 0 1 97920
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_176_197
timestamp 1636968456
transform 1 0 19228 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_209
timestamp 1636968456
transform 1 0 20332 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_221
timestamp 1636968456
transform 1 0 21436 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_233
timestamp 1636968456
transform 1 0 22540 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_176_245
timestamp 1
transform 1 0 23644 0 1 97920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_176_251
timestamp 1
transform 1 0 24196 0 1 97920
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_176_253
timestamp 1636968456
transform 1 0 24380 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_265
timestamp 1636968456
transform 1 0 25484 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_277
timestamp 1636968456
transform 1 0 26588 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_289
timestamp 1636968456
transform 1 0 27692 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_176_301
timestamp 1
transform 1 0 28796 0 1 97920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_176_307
timestamp 1
transform 1 0 29348 0 1 97920
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_176_309
timestamp 1636968456
transform 1 0 29532 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_321
timestamp 1636968456
transform 1 0 30636 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_333
timestamp 1636968456
transform 1 0 31740 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_345
timestamp 1636968456
transform 1 0 32844 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_176_357
timestamp 1
transform 1 0 33948 0 1 97920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_176_363
timestamp 1
transform 1 0 34500 0 1 97920
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_176_365
timestamp 1636968456
transform 1 0 34684 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_377
timestamp 1636968456
transform 1 0 35788 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_389
timestamp 1636968456
transform 1 0 36892 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_401
timestamp 1636968456
transform 1 0 37996 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_176_413
timestamp 1
transform 1 0 39100 0 1 97920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_176_419
timestamp 1
transform 1 0 39652 0 1 97920
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_176_421
timestamp 1636968456
transform 1 0 39836 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_433
timestamp 1636968456
transform 1 0 40940 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_445
timestamp 1636968456
transform 1 0 42044 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_457
timestamp 1636968456
transform 1 0 43148 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_176_469
timestamp 1
transform 1 0 44252 0 1 97920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_176_475
timestamp 1
transform 1 0 44804 0 1 97920
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_176_477
timestamp 1636968456
transform 1 0 44988 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_489
timestamp 1636968456
transform 1 0 46092 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_501
timestamp 1636968456
transform 1 0 47196 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_513
timestamp 1636968456
transform 1 0 48300 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_176_525
timestamp 1
transform 1 0 49404 0 1 97920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_176_531
timestamp 1
transform 1 0 49956 0 1 97920
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_176_533
timestamp 1636968456
transform 1 0 50140 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_545
timestamp 1636968456
transform 1 0 51244 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_557
timestamp 1636968456
transform 1 0 52348 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_569
timestamp 1636968456
transform 1 0 53452 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_176_581
timestamp 1
transform 1 0 54556 0 1 97920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_176_587
timestamp 1
transform 1 0 55108 0 1 97920
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_176_589
timestamp 1636968456
transform 1 0 55292 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_601
timestamp 1636968456
transform 1 0 56396 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_613
timestamp 1636968456
transform 1 0 57500 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_625
timestamp 1636968456
transform 1 0 58604 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_176_637
timestamp 1
transform 1 0 59708 0 1 97920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_176_643
timestamp 1
transform 1 0 60260 0 1 97920
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_176_645
timestamp 1636968456
transform 1 0 60444 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_657
timestamp 1636968456
transform 1 0 61548 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_669
timestamp 1636968456
transform 1 0 62652 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_681
timestamp 1636968456
transform 1 0 63756 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_176_693
timestamp 1
transform 1 0 64860 0 1 97920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_176_699
timestamp 1
transform 1 0 65412 0 1 97920
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_176_701
timestamp 1636968456
transform 1 0 65596 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_713
timestamp 1636968456
transform 1 0 66700 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_725
timestamp 1636968456
transform 1 0 67804 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_737
timestamp 1636968456
transform 1 0 68908 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_176_749
timestamp 1
transform 1 0 70012 0 1 97920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_176_755
timestamp 1
transform 1 0 70564 0 1 97920
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_176_757
timestamp 1636968456
transform 1 0 70748 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_769
timestamp 1636968456
transform 1 0 71852 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_781
timestamp 1636968456
transform 1 0 72956 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_793
timestamp 1636968456
transform 1 0 74060 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_176_805
timestamp 1
transform 1 0 75164 0 1 97920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_176_811
timestamp 1
transform 1 0 75716 0 1 97920
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_176_813
timestamp 1636968456
transform 1 0 75900 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_825
timestamp 1636968456
transform 1 0 77004 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_837
timestamp 1636968456
transform 1 0 78108 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_849
timestamp 1636968456
transform 1 0 79212 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_176_861
timestamp 1
transform 1 0 80316 0 1 97920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_176_867
timestamp 1
transform 1 0 80868 0 1 97920
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_176_869
timestamp 1636968456
transform 1 0 81052 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_881
timestamp 1636968456
transform 1 0 82156 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_893
timestamp 1636968456
transform 1 0 83260 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_905
timestamp 1636968456
transform 1 0 84364 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_176_917
timestamp 1
transform 1 0 85468 0 1 97920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_176_923
timestamp 1
transform 1 0 86020 0 1 97920
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_176_925
timestamp 1636968456
transform 1 0 86204 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_937
timestamp 1636968456
transform 1 0 87308 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_949
timestamp 1636968456
transform 1 0 88412 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_961
timestamp 1636968456
transform 1 0 89516 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_176_973
timestamp 1
transform 1 0 90620 0 1 97920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_176_979
timestamp 1
transform 1 0 91172 0 1 97920
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_176_981
timestamp 1636968456
transform 1 0 91356 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_993
timestamp 1636968456
transform 1 0 92460 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_1005
timestamp 1636968456
transform 1 0 93564 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_1017
timestamp 1636968456
transform 1 0 94668 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_176_1029
timestamp 1
transform 1 0 95772 0 1 97920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_176_1035
timestamp 1
transform 1 0 96324 0 1 97920
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_176_1037
timestamp 1636968456
transform 1 0 96508 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_1049
timestamp 1636968456
transform 1 0 97612 0 1 97920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_176_1061
timestamp 1636968456
transform 1 0 98716 0 1 97920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_176_1073
timestamp 1
transform 1 0 99820 0 1 97920
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_177_3
timestamp 1636968456
transform 1 0 1380 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_15
timestamp 1636968456
transform 1 0 2484 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_27
timestamp 1636968456
transform 1 0 3588 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_39
timestamp 1636968456
transform 1 0 4692 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_177_51
timestamp 1
transform 1 0 5796 0 -1 99008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_177_55
timestamp 1
transform 1 0 6164 0 -1 99008
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_177_57
timestamp 1636968456
transform 1 0 6348 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_69
timestamp 1636968456
transform 1 0 7452 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_81
timestamp 1636968456
transform 1 0 8556 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_93
timestamp 1636968456
transform 1 0 9660 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_177_105
timestamp 1
transform 1 0 10764 0 -1 99008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_177_111
timestamp 1
transform 1 0 11316 0 -1 99008
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_177_113
timestamp 1636968456
transform 1 0 11500 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_125
timestamp 1636968456
transform 1 0 12604 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_137
timestamp 1636968456
transform 1 0 13708 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_149
timestamp 1636968456
transform 1 0 14812 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_177_161
timestamp 1
transform 1 0 15916 0 -1 99008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_177_167
timestamp 1
transform 1 0 16468 0 -1 99008
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_177_169
timestamp 1636968456
transform 1 0 16652 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_181
timestamp 1636968456
transform 1 0 17756 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_193
timestamp 1636968456
transform 1 0 18860 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_205
timestamp 1636968456
transform 1 0 19964 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_177_217
timestamp 1
transform 1 0 21068 0 -1 99008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_177_223
timestamp 1
transform 1 0 21620 0 -1 99008
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_177_225
timestamp 1636968456
transform 1 0 21804 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_237
timestamp 1636968456
transform 1 0 22908 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_249
timestamp 1636968456
transform 1 0 24012 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_261
timestamp 1636968456
transform 1 0 25116 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_177_273
timestamp 1
transform 1 0 26220 0 -1 99008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_177_279
timestamp 1
transform 1 0 26772 0 -1 99008
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_177_281
timestamp 1636968456
transform 1 0 26956 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_293
timestamp 1636968456
transform 1 0 28060 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_305
timestamp 1636968456
transform 1 0 29164 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_317
timestamp 1636968456
transform 1 0 30268 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_177_329
timestamp 1
transform 1 0 31372 0 -1 99008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_177_335
timestamp 1
transform 1 0 31924 0 -1 99008
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_177_337
timestamp 1636968456
transform 1 0 32108 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_349
timestamp 1636968456
transform 1 0 33212 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_361
timestamp 1636968456
transform 1 0 34316 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_373
timestamp 1636968456
transform 1 0 35420 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_177_385
timestamp 1
transform 1 0 36524 0 -1 99008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_177_391
timestamp 1
transform 1 0 37076 0 -1 99008
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_177_393
timestamp 1636968456
transform 1 0 37260 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_405
timestamp 1636968456
transform 1 0 38364 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_417
timestamp 1636968456
transform 1 0 39468 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_429
timestamp 1636968456
transform 1 0 40572 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_177_441
timestamp 1
transform 1 0 41676 0 -1 99008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_177_447
timestamp 1
transform 1 0 42228 0 -1 99008
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_177_449
timestamp 1636968456
transform 1 0 42412 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_461
timestamp 1636968456
transform 1 0 43516 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_473
timestamp 1636968456
transform 1 0 44620 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_485
timestamp 1636968456
transform 1 0 45724 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_177_497
timestamp 1
transform 1 0 46828 0 -1 99008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_177_503
timestamp 1
transform 1 0 47380 0 -1 99008
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_177_505
timestamp 1636968456
transform 1 0 47564 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_517
timestamp 1636968456
transform 1 0 48668 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_529
timestamp 1636968456
transform 1 0 49772 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_541
timestamp 1636968456
transform 1 0 50876 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_177_553
timestamp 1
transform 1 0 51980 0 -1 99008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_177_559
timestamp 1
transform 1 0 52532 0 -1 99008
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_177_561
timestamp 1636968456
transform 1 0 52716 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_573
timestamp 1636968456
transform 1 0 53820 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_585
timestamp 1636968456
transform 1 0 54924 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_597
timestamp 1636968456
transform 1 0 56028 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_177_609
timestamp 1
transform 1 0 57132 0 -1 99008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_177_615
timestamp 1
transform 1 0 57684 0 -1 99008
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_177_617
timestamp 1636968456
transform 1 0 57868 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_629
timestamp 1636968456
transform 1 0 58972 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_641
timestamp 1636968456
transform 1 0 60076 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_653
timestamp 1636968456
transform 1 0 61180 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_177_665
timestamp 1
transform 1 0 62284 0 -1 99008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_177_671
timestamp 1
transform 1 0 62836 0 -1 99008
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_177_673
timestamp 1636968456
transform 1 0 63020 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_685
timestamp 1636968456
transform 1 0 64124 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_697
timestamp 1636968456
transform 1 0 65228 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_709
timestamp 1636968456
transform 1 0 66332 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_177_721
timestamp 1
transform 1 0 67436 0 -1 99008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_177_727
timestamp 1
transform 1 0 67988 0 -1 99008
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_177_729
timestamp 1636968456
transform 1 0 68172 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_741
timestamp 1636968456
transform 1 0 69276 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_753
timestamp 1636968456
transform 1 0 70380 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_765
timestamp 1636968456
transform 1 0 71484 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_177_777
timestamp 1
transform 1 0 72588 0 -1 99008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_177_783
timestamp 1
transform 1 0 73140 0 -1 99008
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_177_785
timestamp 1636968456
transform 1 0 73324 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_797
timestamp 1636968456
transform 1 0 74428 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_809
timestamp 1636968456
transform 1 0 75532 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_821
timestamp 1636968456
transform 1 0 76636 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_177_833
timestamp 1
transform 1 0 77740 0 -1 99008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_177_839
timestamp 1
transform 1 0 78292 0 -1 99008
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_177_841
timestamp 1636968456
transform 1 0 78476 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_853
timestamp 1636968456
transform 1 0 79580 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_865
timestamp 1636968456
transform 1 0 80684 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_877
timestamp 1636968456
transform 1 0 81788 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_177_889
timestamp 1
transform 1 0 82892 0 -1 99008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_177_895
timestamp 1
transform 1 0 83444 0 -1 99008
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_177_897
timestamp 1636968456
transform 1 0 83628 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_909
timestamp 1636968456
transform 1 0 84732 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_921
timestamp 1636968456
transform 1 0 85836 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_933
timestamp 1636968456
transform 1 0 86940 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_177_945
timestamp 1
transform 1 0 88044 0 -1 99008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_177_951
timestamp 1
transform 1 0 88596 0 -1 99008
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_177_953
timestamp 1636968456
transform 1 0 88780 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_965
timestamp 1636968456
transform 1 0 89884 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_977
timestamp 1636968456
transform 1 0 90988 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_989
timestamp 1636968456
transform 1 0 92092 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_177_1001
timestamp 1
transform 1 0 93196 0 -1 99008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_177_1007
timestamp 1
transform 1 0 93748 0 -1 99008
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_177_1009
timestamp 1636968456
transform 1 0 93932 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_1021
timestamp 1636968456
transform 1 0 95036 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_1033
timestamp 1636968456
transform 1 0 96140 0 -1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_177_1045
timestamp 1636968456
transform 1 0 97244 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_177_1057
timestamp 1
transform 1 0 98348 0 -1 99008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_177_1063
timestamp 1
transform 1 0 98900 0 -1 99008
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_177_1065
timestamp 1636968456
transform 1 0 99084 0 -1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_177_1077
timestamp 1
transform 1 0 100188 0 -1 99008
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_178_3
timestamp 1636968456
transform 1 0 1380 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_15
timestamp 1636968456
transform 1 0 2484 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_178_27
timestamp 1
transform 1 0 3588 0 1 99008
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_178_29
timestamp 1636968456
transform 1 0 3772 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_41
timestamp 1636968456
transform 1 0 4876 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_53
timestamp 1636968456
transform 1 0 5980 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_65
timestamp 1636968456
transform 1 0 7084 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_178_77
timestamp 1
transform 1 0 8188 0 1 99008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_178_83
timestamp 1
transform 1 0 8740 0 1 99008
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_178_85
timestamp 1636968456
transform 1 0 8924 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_97
timestamp 1636968456
transform 1 0 10028 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_109
timestamp 1636968456
transform 1 0 11132 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_121
timestamp 1636968456
transform 1 0 12236 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_178_133
timestamp 1
transform 1 0 13340 0 1 99008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_178_139
timestamp 1
transform 1 0 13892 0 1 99008
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_178_141
timestamp 1636968456
transform 1 0 14076 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_153
timestamp 1636968456
transform 1 0 15180 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_165
timestamp 1636968456
transform 1 0 16284 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_177
timestamp 1636968456
transform 1 0 17388 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_178_189
timestamp 1
transform 1 0 18492 0 1 99008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_178_195
timestamp 1
transform 1 0 19044 0 1 99008
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_178_197
timestamp 1636968456
transform 1 0 19228 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_209
timestamp 1636968456
transform 1 0 20332 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_221
timestamp 1636968456
transform 1 0 21436 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_233
timestamp 1636968456
transform 1 0 22540 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_178_245
timestamp 1
transform 1 0 23644 0 1 99008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_178_251
timestamp 1
transform 1 0 24196 0 1 99008
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_178_253
timestamp 1636968456
transform 1 0 24380 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_265
timestamp 1636968456
transform 1 0 25484 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_277
timestamp 1636968456
transform 1 0 26588 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_289
timestamp 1636968456
transform 1 0 27692 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_178_301
timestamp 1
transform 1 0 28796 0 1 99008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_178_307
timestamp 1
transform 1 0 29348 0 1 99008
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_178_309
timestamp 1636968456
transform 1 0 29532 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_321
timestamp 1636968456
transform 1 0 30636 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_333
timestamp 1636968456
transform 1 0 31740 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_345
timestamp 1636968456
transform 1 0 32844 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_178_357
timestamp 1
transform 1 0 33948 0 1 99008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_178_363
timestamp 1
transform 1 0 34500 0 1 99008
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_178_365
timestamp 1636968456
transform 1 0 34684 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_377
timestamp 1636968456
transform 1 0 35788 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_389
timestamp 1636968456
transform 1 0 36892 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_401
timestamp 1636968456
transform 1 0 37996 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_178_413
timestamp 1
transform 1 0 39100 0 1 99008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_178_419
timestamp 1
transform 1 0 39652 0 1 99008
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_178_421
timestamp 1636968456
transform 1 0 39836 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_433
timestamp 1636968456
transform 1 0 40940 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_445
timestamp 1636968456
transform 1 0 42044 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_457
timestamp 1636968456
transform 1 0 43148 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_178_469
timestamp 1
transform 1 0 44252 0 1 99008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_178_475
timestamp 1
transform 1 0 44804 0 1 99008
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_178_477
timestamp 1636968456
transform 1 0 44988 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_489
timestamp 1636968456
transform 1 0 46092 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_501
timestamp 1636968456
transform 1 0 47196 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_513
timestamp 1636968456
transform 1 0 48300 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_178_525
timestamp 1
transform 1 0 49404 0 1 99008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_178_531
timestamp 1
transform 1 0 49956 0 1 99008
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_178_533
timestamp 1636968456
transform 1 0 50140 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_545
timestamp 1636968456
transform 1 0 51244 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_557
timestamp 1636968456
transform 1 0 52348 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_569
timestamp 1636968456
transform 1 0 53452 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_178_581
timestamp 1
transform 1 0 54556 0 1 99008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_178_587
timestamp 1
transform 1 0 55108 0 1 99008
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_178_589
timestamp 1636968456
transform 1 0 55292 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_601
timestamp 1636968456
transform 1 0 56396 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_613
timestamp 1636968456
transform 1 0 57500 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_625
timestamp 1636968456
transform 1 0 58604 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_178_637
timestamp 1
transform 1 0 59708 0 1 99008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_178_643
timestamp 1
transform 1 0 60260 0 1 99008
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_178_645
timestamp 1636968456
transform 1 0 60444 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_657
timestamp 1636968456
transform 1 0 61548 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_669
timestamp 1636968456
transform 1 0 62652 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_681
timestamp 1636968456
transform 1 0 63756 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_178_693
timestamp 1
transform 1 0 64860 0 1 99008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_178_699
timestamp 1
transform 1 0 65412 0 1 99008
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_178_701
timestamp 1636968456
transform 1 0 65596 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_713
timestamp 1636968456
transform 1 0 66700 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_725
timestamp 1636968456
transform 1 0 67804 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_737
timestamp 1636968456
transform 1 0 68908 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_178_749
timestamp 1
transform 1 0 70012 0 1 99008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_178_755
timestamp 1
transform 1 0 70564 0 1 99008
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_178_757
timestamp 1636968456
transform 1 0 70748 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_769
timestamp 1636968456
transform 1 0 71852 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_781
timestamp 1636968456
transform 1 0 72956 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_793
timestamp 1636968456
transform 1 0 74060 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_178_805
timestamp 1
transform 1 0 75164 0 1 99008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_178_811
timestamp 1
transform 1 0 75716 0 1 99008
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_178_813
timestamp 1636968456
transform 1 0 75900 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_825
timestamp 1636968456
transform 1 0 77004 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_837
timestamp 1636968456
transform 1 0 78108 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_849
timestamp 1636968456
transform 1 0 79212 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_178_861
timestamp 1
transform 1 0 80316 0 1 99008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_178_867
timestamp 1
transform 1 0 80868 0 1 99008
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_178_869
timestamp 1636968456
transform 1 0 81052 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_881
timestamp 1636968456
transform 1 0 82156 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_893
timestamp 1636968456
transform 1 0 83260 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_905
timestamp 1636968456
transform 1 0 84364 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_178_917
timestamp 1
transform 1 0 85468 0 1 99008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_178_923
timestamp 1
transform 1 0 86020 0 1 99008
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_178_925
timestamp 1636968456
transform 1 0 86204 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_937
timestamp 1636968456
transform 1 0 87308 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_949
timestamp 1636968456
transform 1 0 88412 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_961
timestamp 1636968456
transform 1 0 89516 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_178_973
timestamp 1
transform 1 0 90620 0 1 99008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_178_979
timestamp 1
transform 1 0 91172 0 1 99008
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_178_981
timestamp 1636968456
transform 1 0 91356 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_993
timestamp 1636968456
transform 1 0 92460 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_1005
timestamp 1636968456
transform 1 0 93564 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_1017
timestamp 1636968456
transform 1 0 94668 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_178_1029
timestamp 1
transform 1 0 95772 0 1 99008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_178_1035
timestamp 1
transform 1 0 96324 0 1 99008
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_178_1037
timestamp 1636968456
transform 1 0 96508 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_1049
timestamp 1636968456
transform 1 0 97612 0 1 99008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_178_1061
timestamp 1636968456
transform 1 0 98716 0 1 99008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_178_1073
timestamp 1
transform 1 0 99820 0 1 99008
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_179_3
timestamp 1636968456
transform 1 0 1380 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_15
timestamp 1636968456
transform 1 0 2484 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_27
timestamp 1636968456
transform 1 0 3588 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_39
timestamp 1636968456
transform 1 0 4692 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_179_51
timestamp 1
transform 1 0 5796 0 -1 100096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_179_55
timestamp 1
transform 1 0 6164 0 -1 100096
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_179_57
timestamp 1636968456
transform 1 0 6348 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_69
timestamp 1636968456
transform 1 0 7452 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_81
timestamp 1636968456
transform 1 0 8556 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_93
timestamp 1636968456
transform 1 0 9660 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_179_105
timestamp 1
transform 1 0 10764 0 -1 100096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_179_111
timestamp 1
transform 1 0 11316 0 -1 100096
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_179_113
timestamp 1636968456
transform 1 0 11500 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_125
timestamp 1636968456
transform 1 0 12604 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_137
timestamp 1636968456
transform 1 0 13708 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_149
timestamp 1636968456
transform 1 0 14812 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_179_161
timestamp 1
transform 1 0 15916 0 -1 100096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_179_167
timestamp 1
transform 1 0 16468 0 -1 100096
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_179_169
timestamp 1636968456
transform 1 0 16652 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_181
timestamp 1636968456
transform 1 0 17756 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_193
timestamp 1636968456
transform 1 0 18860 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_205
timestamp 1636968456
transform 1 0 19964 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_179_217
timestamp 1
transform 1 0 21068 0 -1 100096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_179_223
timestamp 1
transform 1 0 21620 0 -1 100096
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_179_225
timestamp 1636968456
transform 1 0 21804 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_237
timestamp 1636968456
transform 1 0 22908 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_249
timestamp 1636968456
transform 1 0 24012 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_261
timestamp 1636968456
transform 1 0 25116 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_179_273
timestamp 1
transform 1 0 26220 0 -1 100096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_179_279
timestamp 1
transform 1 0 26772 0 -1 100096
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_179_281
timestamp 1636968456
transform 1 0 26956 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_293
timestamp 1636968456
transform 1 0 28060 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_305
timestamp 1636968456
transform 1 0 29164 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_317
timestamp 1636968456
transform 1 0 30268 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_179_329
timestamp 1
transform 1 0 31372 0 -1 100096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_179_335
timestamp 1
transform 1 0 31924 0 -1 100096
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_179_337
timestamp 1636968456
transform 1 0 32108 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_349
timestamp 1636968456
transform 1 0 33212 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_361
timestamp 1636968456
transform 1 0 34316 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_373
timestamp 1636968456
transform 1 0 35420 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_179_385
timestamp 1
transform 1 0 36524 0 -1 100096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_179_391
timestamp 1
transform 1 0 37076 0 -1 100096
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_179_393
timestamp 1636968456
transform 1 0 37260 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_405
timestamp 1636968456
transform 1 0 38364 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_417
timestamp 1636968456
transform 1 0 39468 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_429
timestamp 1636968456
transform 1 0 40572 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_179_441
timestamp 1
transform 1 0 41676 0 -1 100096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_179_447
timestamp 1
transform 1 0 42228 0 -1 100096
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_179_449
timestamp 1636968456
transform 1 0 42412 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_461
timestamp 1636968456
transform 1 0 43516 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_473
timestamp 1636968456
transform 1 0 44620 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_485
timestamp 1636968456
transform 1 0 45724 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_179_497
timestamp 1
transform 1 0 46828 0 -1 100096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_179_503
timestamp 1
transform 1 0 47380 0 -1 100096
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_179_505
timestamp 1636968456
transform 1 0 47564 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_517
timestamp 1636968456
transform 1 0 48668 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_529
timestamp 1636968456
transform 1 0 49772 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_541
timestamp 1636968456
transform 1 0 50876 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_179_553
timestamp 1
transform 1 0 51980 0 -1 100096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_179_559
timestamp 1
transform 1 0 52532 0 -1 100096
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_179_561
timestamp 1636968456
transform 1 0 52716 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_573
timestamp 1636968456
transform 1 0 53820 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_585
timestamp 1636968456
transform 1 0 54924 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_597
timestamp 1636968456
transform 1 0 56028 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_179_609
timestamp 1
transform 1 0 57132 0 -1 100096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_179_615
timestamp 1
transform 1 0 57684 0 -1 100096
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_179_617
timestamp 1636968456
transform 1 0 57868 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_629
timestamp 1636968456
transform 1 0 58972 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_641
timestamp 1636968456
transform 1 0 60076 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_653
timestamp 1636968456
transform 1 0 61180 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_179_665
timestamp 1
transform 1 0 62284 0 -1 100096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_179_671
timestamp 1
transform 1 0 62836 0 -1 100096
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_179_673
timestamp 1636968456
transform 1 0 63020 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_685
timestamp 1636968456
transform 1 0 64124 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_697
timestamp 1636968456
transform 1 0 65228 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_709
timestamp 1636968456
transform 1 0 66332 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_179_721
timestamp 1
transform 1 0 67436 0 -1 100096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_179_727
timestamp 1
transform 1 0 67988 0 -1 100096
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_179_729
timestamp 1636968456
transform 1 0 68172 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_741
timestamp 1636968456
transform 1 0 69276 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_753
timestamp 1636968456
transform 1 0 70380 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_765
timestamp 1636968456
transform 1 0 71484 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_179_777
timestamp 1
transform 1 0 72588 0 -1 100096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_179_783
timestamp 1
transform 1 0 73140 0 -1 100096
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_179_785
timestamp 1636968456
transform 1 0 73324 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_797
timestamp 1636968456
transform 1 0 74428 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_809
timestamp 1636968456
transform 1 0 75532 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_821
timestamp 1636968456
transform 1 0 76636 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_179_833
timestamp 1
transform 1 0 77740 0 -1 100096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_179_839
timestamp 1
transform 1 0 78292 0 -1 100096
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_179_841
timestamp 1636968456
transform 1 0 78476 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_853
timestamp 1636968456
transform 1 0 79580 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_865
timestamp 1636968456
transform 1 0 80684 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_877
timestamp 1636968456
transform 1 0 81788 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_179_889
timestamp 1
transform 1 0 82892 0 -1 100096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_179_895
timestamp 1
transform 1 0 83444 0 -1 100096
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_179_897
timestamp 1636968456
transform 1 0 83628 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_909
timestamp 1636968456
transform 1 0 84732 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_921
timestamp 1636968456
transform 1 0 85836 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_933
timestamp 1636968456
transform 1 0 86940 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_179_945
timestamp 1
transform 1 0 88044 0 -1 100096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_179_951
timestamp 1
transform 1 0 88596 0 -1 100096
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_179_953
timestamp 1636968456
transform 1 0 88780 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_965
timestamp 1636968456
transform 1 0 89884 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_977
timestamp 1636968456
transform 1 0 90988 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_989
timestamp 1636968456
transform 1 0 92092 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_179_1001
timestamp 1
transform 1 0 93196 0 -1 100096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_179_1007
timestamp 1
transform 1 0 93748 0 -1 100096
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_179_1009
timestamp 1636968456
transform 1 0 93932 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_1021
timestamp 1636968456
transform 1 0 95036 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_1033
timestamp 1636968456
transform 1 0 96140 0 -1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_179_1045
timestamp 1636968456
transform 1 0 97244 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_179_1057
timestamp 1
transform 1 0 98348 0 -1 100096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_179_1063
timestamp 1
transform 1 0 98900 0 -1 100096
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_179_1065
timestamp 1636968456
transform 1 0 99084 0 -1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_179_1077
timestamp 1
transform 1 0 100188 0 -1 100096
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_180_3
timestamp 1636968456
transform 1 0 1380 0 1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_180_15
timestamp 1636968456
transform 1 0 2484 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_180_27
timestamp 1
transform 1 0 3588 0 1 100096
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_180_29
timestamp 1636968456
transform 1 0 3772 0 1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_180_41
timestamp 1636968456
transform 1 0 4876 0 1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_180_53
timestamp 1636968456
transform 1 0 5980 0 1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_180_65
timestamp 1636968456
transform 1 0 7084 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_180_77
timestamp 1
transform 1 0 8188 0 1 100096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_180_83
timestamp 1
transform 1 0 8740 0 1 100096
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_180_85
timestamp 1636968456
transform 1 0 8924 0 1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_180_97
timestamp 1636968456
transform 1 0 10028 0 1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_180_109
timestamp 1636968456
transform 1 0 11132 0 1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_180_121
timestamp 1636968456
transform 1 0 12236 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_180_133
timestamp 1
transform 1 0 13340 0 1 100096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_180_139
timestamp 1
transform 1 0 13892 0 1 100096
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_180_141
timestamp 1636968456
transform 1 0 14076 0 1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_180_153
timestamp 1636968456
transform 1 0 15180 0 1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_180_165
timestamp 1636968456
transform 1 0 16284 0 1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_180_177
timestamp 1636968456
transform 1 0 17388 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_180_189
timestamp 1
transform 1 0 18492 0 1 100096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_180_195
timestamp 1
transform 1 0 19044 0 1 100096
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_180_197
timestamp 1636968456
transform 1 0 19228 0 1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_180_209
timestamp 1636968456
transform 1 0 20332 0 1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_180_221
timestamp 1636968456
transform 1 0 21436 0 1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_180_233
timestamp 1636968456
transform 1 0 22540 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_180_245
timestamp 1
transform 1 0 23644 0 1 100096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_180_251
timestamp 1
transform 1 0 24196 0 1 100096
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_180_253
timestamp 1636968456
transform 1 0 24380 0 1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_180_265
timestamp 1636968456
transform 1 0 25484 0 1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_180_277
timestamp 1636968456
transform 1 0 26588 0 1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_180_289
timestamp 1636968456
transform 1 0 27692 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_180_301
timestamp 1
transform 1 0 28796 0 1 100096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_180_307
timestamp 1
transform 1 0 29348 0 1 100096
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_180_309
timestamp 1636968456
transform 1 0 29532 0 1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_180_321
timestamp 1636968456
transform 1 0 30636 0 1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_180_333
timestamp 1636968456
transform 1 0 31740 0 1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_180_345
timestamp 1636968456
transform 1 0 32844 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_180_357
timestamp 1
transform 1 0 33948 0 1 100096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_180_363
timestamp 1
transform 1 0 34500 0 1 100096
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_180_365
timestamp 1636968456
transform 1 0 34684 0 1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_180_377
timestamp 1636968456
transform 1 0 35788 0 1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_180_389
timestamp 1636968456
transform 1 0 36892 0 1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_180_401
timestamp 1636968456
transform 1 0 37996 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_180_413
timestamp 1
transform 1 0 39100 0 1 100096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_180_419
timestamp 1
transform 1 0 39652 0 1 100096
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_180_421
timestamp 1636968456
transform 1 0 39836 0 1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_180_433
timestamp 1636968456
transform 1 0 40940 0 1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_180_445
timestamp 1636968456
transform 1 0 42044 0 1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_180_457
timestamp 1636968456
transform 1 0 43148 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_180_469
timestamp 1
transform 1 0 44252 0 1 100096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_180_475
timestamp 1
transform 1 0 44804 0 1 100096
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_180_477
timestamp 1636968456
transform 1 0 44988 0 1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_180_489
timestamp 1636968456
transform 1 0 46092 0 1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_180_501
timestamp 1636968456
transform 1 0 47196 0 1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_180_513
timestamp 1636968456
transform 1 0 48300 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_180_525
timestamp 1
transform 1 0 49404 0 1 100096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_180_531
timestamp 1
transform 1 0 49956 0 1 100096
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_180_533
timestamp 1636968456
transform 1 0 50140 0 1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_180_545
timestamp 1636968456
transform 1 0 51244 0 1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_180_557
timestamp 1636968456
transform 1 0 52348 0 1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_180_569
timestamp 1636968456
transform 1 0 53452 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_180_581
timestamp 1
transform 1 0 54556 0 1 100096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_180_587
timestamp 1
transform 1 0 55108 0 1 100096
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_180_589
timestamp 1636968456
transform 1 0 55292 0 1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_180_601
timestamp 1636968456
transform 1 0 56396 0 1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_180_613
timestamp 1636968456
transform 1 0 57500 0 1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_180_625
timestamp 1636968456
transform 1 0 58604 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_180_637
timestamp 1
transform 1 0 59708 0 1 100096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_180_643
timestamp 1
transform 1 0 60260 0 1 100096
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_180_645
timestamp 1636968456
transform 1 0 60444 0 1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_180_657
timestamp 1636968456
transform 1 0 61548 0 1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_180_669
timestamp 1636968456
transform 1 0 62652 0 1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_180_681
timestamp 1636968456
transform 1 0 63756 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_180_693
timestamp 1
transform 1 0 64860 0 1 100096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_180_699
timestamp 1
transform 1 0 65412 0 1 100096
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_180_701
timestamp 1636968456
transform 1 0 65596 0 1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_180_713
timestamp 1636968456
transform 1 0 66700 0 1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_180_725
timestamp 1636968456
transform 1 0 67804 0 1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_180_737
timestamp 1636968456
transform 1 0 68908 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_180_749
timestamp 1
transform 1 0 70012 0 1 100096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_180_755
timestamp 1
transform 1 0 70564 0 1 100096
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_180_757
timestamp 1636968456
transform 1 0 70748 0 1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_180_769
timestamp 1636968456
transform 1 0 71852 0 1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_180_781
timestamp 1636968456
transform 1 0 72956 0 1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_180_793
timestamp 1636968456
transform 1 0 74060 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_180_805
timestamp 1
transform 1 0 75164 0 1 100096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_180_811
timestamp 1
transform 1 0 75716 0 1 100096
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_180_813
timestamp 1636968456
transform 1 0 75900 0 1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_180_825
timestamp 1636968456
transform 1 0 77004 0 1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_180_837
timestamp 1636968456
transform 1 0 78108 0 1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_180_849
timestamp 1636968456
transform 1 0 79212 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_180_861
timestamp 1
transform 1 0 80316 0 1 100096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_180_867
timestamp 1
transform 1 0 80868 0 1 100096
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_180_869
timestamp 1636968456
transform 1 0 81052 0 1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_180_881
timestamp 1636968456
transform 1 0 82156 0 1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_180_893
timestamp 1636968456
transform 1 0 83260 0 1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_180_905
timestamp 1636968456
transform 1 0 84364 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_180_917
timestamp 1
transform 1 0 85468 0 1 100096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_180_923
timestamp 1
transform 1 0 86020 0 1 100096
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_180_925
timestamp 1636968456
transform 1 0 86204 0 1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_180_937
timestamp 1636968456
transform 1 0 87308 0 1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_180_949
timestamp 1636968456
transform 1 0 88412 0 1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_180_961
timestamp 1636968456
transform 1 0 89516 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_180_973
timestamp 1
transform 1 0 90620 0 1 100096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_180_979
timestamp 1
transform 1 0 91172 0 1 100096
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_180_981
timestamp 1636968456
transform 1 0 91356 0 1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_180_993
timestamp 1636968456
transform 1 0 92460 0 1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_180_1005
timestamp 1636968456
transform 1 0 93564 0 1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_180_1017
timestamp 1636968456
transform 1 0 94668 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_180_1029
timestamp 1
transform 1 0 95772 0 1 100096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_180_1035
timestamp 1
transform 1 0 96324 0 1 100096
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_180_1037
timestamp 1636968456
transform 1 0 96508 0 1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_180_1049
timestamp 1636968456
transform 1 0 97612 0 1 100096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_180_1061
timestamp 1636968456
transform 1 0 98716 0 1 100096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_180_1073
timestamp 1
transform 1 0 99820 0 1 100096
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_181_3
timestamp 1636968456
transform 1 0 1380 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_15
timestamp 1636968456
transform 1 0 2484 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_27
timestamp 1636968456
transform 1 0 3588 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_39
timestamp 1636968456
transform 1 0 4692 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_181_51
timestamp 1
transform 1 0 5796 0 -1 101184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_181_55
timestamp 1
transform 1 0 6164 0 -1 101184
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_181_57
timestamp 1636968456
transform 1 0 6348 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_69
timestamp 1636968456
transform 1 0 7452 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_81
timestamp 1636968456
transform 1 0 8556 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_93
timestamp 1636968456
transform 1 0 9660 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_181_105
timestamp 1
transform 1 0 10764 0 -1 101184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_181_111
timestamp 1
transform 1 0 11316 0 -1 101184
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_181_113
timestamp 1636968456
transform 1 0 11500 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_125
timestamp 1636968456
transform 1 0 12604 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_137
timestamp 1636968456
transform 1 0 13708 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_149
timestamp 1636968456
transform 1 0 14812 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_181_161
timestamp 1
transform 1 0 15916 0 -1 101184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_181_167
timestamp 1
transform 1 0 16468 0 -1 101184
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_181_169
timestamp 1636968456
transform 1 0 16652 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_181
timestamp 1636968456
transform 1 0 17756 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_193
timestamp 1636968456
transform 1 0 18860 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_205
timestamp 1636968456
transform 1 0 19964 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_181_217
timestamp 1
transform 1 0 21068 0 -1 101184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_181_223
timestamp 1
transform 1 0 21620 0 -1 101184
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_181_225
timestamp 1636968456
transform 1 0 21804 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_237
timestamp 1636968456
transform 1 0 22908 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_249
timestamp 1636968456
transform 1 0 24012 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_261
timestamp 1636968456
transform 1 0 25116 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_181_273
timestamp 1
transform 1 0 26220 0 -1 101184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_181_279
timestamp 1
transform 1 0 26772 0 -1 101184
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_181_281
timestamp 1636968456
transform 1 0 26956 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_293
timestamp 1636968456
transform 1 0 28060 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_305
timestamp 1636968456
transform 1 0 29164 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_317
timestamp 1636968456
transform 1 0 30268 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_181_329
timestamp 1
transform 1 0 31372 0 -1 101184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_181_335
timestamp 1
transform 1 0 31924 0 -1 101184
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_181_337
timestamp 1636968456
transform 1 0 32108 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_349
timestamp 1636968456
transform 1 0 33212 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_361
timestamp 1636968456
transform 1 0 34316 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_373
timestamp 1636968456
transform 1 0 35420 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_181_385
timestamp 1
transform 1 0 36524 0 -1 101184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_181_391
timestamp 1
transform 1 0 37076 0 -1 101184
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_181_393
timestamp 1636968456
transform 1 0 37260 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_405
timestamp 1636968456
transform 1 0 38364 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_417
timestamp 1636968456
transform 1 0 39468 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_429
timestamp 1636968456
transform 1 0 40572 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_181_441
timestamp 1
transform 1 0 41676 0 -1 101184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_181_447
timestamp 1
transform 1 0 42228 0 -1 101184
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_181_449
timestamp 1636968456
transform 1 0 42412 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_461
timestamp 1636968456
transform 1 0 43516 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_473
timestamp 1636968456
transform 1 0 44620 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_485
timestamp 1636968456
transform 1 0 45724 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_181_497
timestamp 1
transform 1 0 46828 0 -1 101184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_181_503
timestamp 1
transform 1 0 47380 0 -1 101184
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_181_505
timestamp 1636968456
transform 1 0 47564 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_517
timestamp 1636968456
transform 1 0 48668 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_529
timestamp 1636968456
transform 1 0 49772 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_541
timestamp 1636968456
transform 1 0 50876 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_181_553
timestamp 1
transform 1 0 51980 0 -1 101184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_181_559
timestamp 1
transform 1 0 52532 0 -1 101184
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_181_561
timestamp 1636968456
transform 1 0 52716 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_573
timestamp 1636968456
transform 1 0 53820 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_585
timestamp 1636968456
transform 1 0 54924 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_597
timestamp 1636968456
transform 1 0 56028 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_181_609
timestamp 1
transform 1 0 57132 0 -1 101184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_181_615
timestamp 1
transform 1 0 57684 0 -1 101184
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_181_617
timestamp 1636968456
transform 1 0 57868 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_629
timestamp 1636968456
transform 1 0 58972 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_641
timestamp 1636968456
transform 1 0 60076 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_653
timestamp 1636968456
transform 1 0 61180 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_181_665
timestamp 1
transform 1 0 62284 0 -1 101184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_181_671
timestamp 1
transform 1 0 62836 0 -1 101184
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_181_673
timestamp 1636968456
transform 1 0 63020 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_685
timestamp 1636968456
transform 1 0 64124 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_697
timestamp 1636968456
transform 1 0 65228 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_709
timestamp 1636968456
transform 1 0 66332 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_181_721
timestamp 1
transform 1 0 67436 0 -1 101184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_181_727
timestamp 1
transform 1 0 67988 0 -1 101184
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_181_729
timestamp 1636968456
transform 1 0 68172 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_741
timestamp 1636968456
transform 1 0 69276 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_753
timestamp 1636968456
transform 1 0 70380 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_765
timestamp 1636968456
transform 1 0 71484 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_181_777
timestamp 1
transform 1 0 72588 0 -1 101184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_181_783
timestamp 1
transform 1 0 73140 0 -1 101184
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_181_785
timestamp 1636968456
transform 1 0 73324 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_797
timestamp 1636968456
transform 1 0 74428 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_809
timestamp 1636968456
transform 1 0 75532 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_821
timestamp 1636968456
transform 1 0 76636 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_181_833
timestamp 1
transform 1 0 77740 0 -1 101184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_181_839
timestamp 1
transform 1 0 78292 0 -1 101184
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_181_841
timestamp 1636968456
transform 1 0 78476 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_853
timestamp 1636968456
transform 1 0 79580 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_865
timestamp 1636968456
transform 1 0 80684 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_877
timestamp 1636968456
transform 1 0 81788 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_181_889
timestamp 1
transform 1 0 82892 0 -1 101184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_181_895
timestamp 1
transform 1 0 83444 0 -1 101184
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_181_897
timestamp 1636968456
transform 1 0 83628 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_909
timestamp 1636968456
transform 1 0 84732 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_921
timestamp 1636968456
transform 1 0 85836 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_933
timestamp 1636968456
transform 1 0 86940 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_181_945
timestamp 1
transform 1 0 88044 0 -1 101184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_181_951
timestamp 1
transform 1 0 88596 0 -1 101184
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_181_953
timestamp 1636968456
transform 1 0 88780 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_965
timestamp 1636968456
transform 1 0 89884 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_977
timestamp 1636968456
transform 1 0 90988 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_989
timestamp 1636968456
transform 1 0 92092 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_181_1001
timestamp 1
transform 1 0 93196 0 -1 101184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_181_1007
timestamp 1
transform 1 0 93748 0 -1 101184
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_181_1009
timestamp 1636968456
transform 1 0 93932 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_1021
timestamp 1636968456
transform 1 0 95036 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_1033
timestamp 1636968456
transform 1 0 96140 0 -1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_181_1045
timestamp 1636968456
transform 1 0 97244 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_181_1057
timestamp 1
transform 1 0 98348 0 -1 101184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_181_1063
timestamp 1
transform 1 0 98900 0 -1 101184
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_181_1065
timestamp 1636968456
transform 1 0 99084 0 -1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_181_1077
timestamp 1
transform 1 0 100188 0 -1 101184
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_182_3
timestamp 1636968456
transform 1 0 1380 0 1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_182_15
timestamp 1636968456
transform 1 0 2484 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_182_27
timestamp 1
transform 1 0 3588 0 1 101184
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_182_29
timestamp 1636968456
transform 1 0 3772 0 1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_182_41
timestamp 1636968456
transform 1 0 4876 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_182_53
timestamp 1
transform 1 0 5980 0 1 101184
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_182_57
timestamp 1636968456
transform 1 0 6348 0 1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_182_69
timestamp 1636968456
transform 1 0 7452 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_182_81
timestamp 1
transform 1 0 8556 0 1 101184
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_182_85
timestamp 1636968456
transform 1 0 8924 0 1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_182_97
timestamp 1636968456
transform 1 0 10028 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_182_109
timestamp 1
transform 1 0 11132 0 1 101184
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_182_113
timestamp 1636968456
transform 1 0 11500 0 1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_182_125
timestamp 1636968456
transform 1 0 12604 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_182_137
timestamp 1
transform 1 0 13708 0 1 101184
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_182_141
timestamp 1636968456
transform 1 0 14076 0 1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_182_153
timestamp 1636968456
transform 1 0 15180 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_182_165
timestamp 1
transform 1 0 16284 0 1 101184
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_182_169
timestamp 1636968456
transform 1 0 16652 0 1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_182_181
timestamp 1636968456
transform 1 0 17756 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_182_193
timestamp 1
transform 1 0 18860 0 1 101184
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_182_197
timestamp 1636968456
transform 1 0 19228 0 1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_182_209
timestamp 1636968456
transform 1 0 20332 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_182_221
timestamp 1
transform 1 0 21436 0 1 101184
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_182_225
timestamp 1636968456
transform 1 0 21804 0 1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_182_237
timestamp 1636968456
transform 1 0 22908 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_182_249
timestamp 1
transform 1 0 24012 0 1 101184
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_182_253
timestamp 1636968456
transform 1 0 24380 0 1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_182_265
timestamp 1636968456
transform 1 0 25484 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_182_277
timestamp 1
transform 1 0 26588 0 1 101184
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_182_281
timestamp 1636968456
transform 1 0 26956 0 1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_182_293
timestamp 1636968456
transform 1 0 28060 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_182_305
timestamp 1
transform 1 0 29164 0 1 101184
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_182_309
timestamp 1636968456
transform 1 0 29532 0 1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_182_321
timestamp 1636968456
transform 1 0 30636 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_182_333
timestamp 1
transform 1 0 31740 0 1 101184
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_182_337
timestamp 1636968456
transform 1 0 32108 0 1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_182_349
timestamp 1636968456
transform 1 0 33212 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_182_361
timestamp 1
transform 1 0 34316 0 1 101184
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_182_365
timestamp 1636968456
transform 1 0 34684 0 1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_182_377
timestamp 1636968456
transform 1 0 35788 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_182_389
timestamp 1
transform 1 0 36892 0 1 101184
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_182_393
timestamp 1636968456
transform 1 0 37260 0 1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_182_405
timestamp 1636968456
transform 1 0 38364 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_182_417
timestamp 1
transform 1 0 39468 0 1 101184
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_182_421
timestamp 1636968456
transform 1 0 39836 0 1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_182_433
timestamp 1636968456
transform 1 0 40940 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_182_445
timestamp 1
transform 1 0 42044 0 1 101184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_182_449
timestamp 1
transform 1 0 42412 0 1 101184
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_182_457
timestamp 1
transform 1 0 43148 0 1 101184
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_182_462
timestamp 1636968456
transform 1 0 43608 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_182_474
timestamp 1
transform 1 0 44712 0 1 101184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_182_477
timestamp 1
transform 1 0 44988 0 1 101184
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_182_483
timestamp 1636968456
transform 1 0 45540 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_182_495
timestamp 1
transform 1 0 46644 0 1 101184
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_182_503
timestamp 1
transform 1 0 47380 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_182_505
timestamp 1
transform 1 0 47564 0 1 101184
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_182_511
timestamp 1636968456
transform 1 0 48116 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_182_523
timestamp 1
transform 1 0 49220 0 1 101184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_182_527
timestamp 1
transform 1 0 49588 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_182_533
timestamp 1
transform 1 0 50140 0 1 101184
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_182_541
timestamp 1
transform 1 0 50876 0 1 101184
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_182_546
timestamp 1636968456
transform 1 0 51336 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_182_558
timestamp 1
transform 1 0 52440 0 1 101184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_182_561
timestamp 1
transform 1 0 52716 0 1 101184
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_182_567
timestamp 1636968456
transform 1 0 53268 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_182_579
timestamp 1
transform 1 0 54372 0 1 101184
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_182_587
timestamp 1
transform 1 0 55108 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_182_589
timestamp 1
transform 1 0 55292 0 1 101184
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_182_595
timestamp 1636968456
transform 1 0 55844 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_182_607
timestamp 1
transform 1 0 56948 0 1 101184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_182_611
timestamp 1
transform 1 0 57316 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_182_617
timestamp 1
transform 1 0 57868 0 1 101184
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_182_625
timestamp 1
transform 1 0 58604 0 1 101184
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_182_630
timestamp 1636968456
transform 1 0 59064 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_182_642
timestamp 1
transform 1 0 60168 0 1 101184
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_182_645
timestamp 1636968456
transform 1 0 60444 0 1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_182_657
timestamp 1636968456
transform 1 0 61548 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_182_669
timestamp 1
transform 1 0 62652 0 1 101184
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_182_673
timestamp 1636968456
transform 1 0 63020 0 1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_182_685
timestamp 1636968456
transform 1 0 64124 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_182_697
timestamp 1
transform 1 0 65228 0 1 101184
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_182_701
timestamp 1636968456
transform 1 0 65596 0 1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_182_713
timestamp 1636968456
transform 1 0 66700 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_182_725
timestamp 1
transform 1 0 67804 0 1 101184
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_182_729
timestamp 1636968456
transform 1 0 68172 0 1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_182_741
timestamp 1636968456
transform 1 0 69276 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_182_753
timestamp 1
transform 1 0 70380 0 1 101184
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_182_757
timestamp 1636968456
transform 1 0 70748 0 1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_182_769
timestamp 1636968456
transform 1 0 71852 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_182_781
timestamp 1
transform 1 0 72956 0 1 101184
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_182_785
timestamp 1636968456
transform 1 0 73324 0 1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_182_797
timestamp 1636968456
transform 1 0 74428 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_182_809
timestamp 1
transform 1 0 75532 0 1 101184
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_182_813
timestamp 1636968456
transform 1 0 75900 0 1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_182_825
timestamp 1636968456
transform 1 0 77004 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_182_837
timestamp 1
transform 1 0 78108 0 1 101184
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_182_841
timestamp 1636968456
transform 1 0 78476 0 1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_182_853
timestamp 1636968456
transform 1 0 79580 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_182_865
timestamp 1
transform 1 0 80684 0 1 101184
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_182_869
timestamp 1636968456
transform 1 0 81052 0 1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_182_881
timestamp 1636968456
transform 1 0 82156 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_182_893
timestamp 1
transform 1 0 83260 0 1 101184
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_182_897
timestamp 1636968456
transform 1 0 83628 0 1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_182_909
timestamp 1636968456
transform 1 0 84732 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_182_921
timestamp 1
transform 1 0 85836 0 1 101184
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_182_925
timestamp 1636968456
transform 1 0 86204 0 1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_182_937
timestamp 1636968456
transform 1 0 87308 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_182_949
timestamp 1
transform 1 0 88412 0 1 101184
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_182_953
timestamp 1636968456
transform 1 0 88780 0 1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_182_965
timestamp 1636968456
transform 1 0 89884 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_182_977
timestamp 1
transform 1 0 90988 0 1 101184
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_182_981
timestamp 1636968456
transform 1 0 91356 0 1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_182_993
timestamp 1636968456
transform 1 0 92460 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_182_1005
timestamp 1
transform 1 0 93564 0 1 101184
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_182_1009
timestamp 1636968456
transform 1 0 93932 0 1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_182_1021
timestamp 1636968456
transform 1 0 95036 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_182_1033
timestamp 1
transform 1 0 96140 0 1 101184
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_182_1037
timestamp 1636968456
transform 1 0 96508 0 1 101184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_182_1049
timestamp 1636968456
transform 1 0 97612 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_182_1061
timestamp 1
transform 1 0 98716 0 1 101184
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_182_1065
timestamp 1636968456
transform 1 0 99084 0 1 101184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_182_1077
timestamp 1
transform 1 0 100188 0 1 101184
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp 1
transform -1 0 99176 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1
transform 1 0 85100 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1
transform 1 0 98716 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1
transform 1 0 86940 0 1 59840
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1
transform 1 0 98808 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1
transform 1 0 100280 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mem_i_21
timestamp 1
transform -1 0 98532 0 -1 54400
box -38 -48 314 592
use ram256x16  mem_i
timestamp 0
transform 1 0 4000 0 1 4000
box 0 0 1 1
use sky130_fd_sc_hd__buf_2  output2
timestamp 1
transform -1 0 1748 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output3
timestamp 1
transform -1 0 59064 0 1 101184
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output4
timestamp 1
transform 1 0 100188 0 -1 63104
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output5
timestamp 1
transform 1 0 100188 0 1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output6
timestamp 1
transform 1 0 100188 0 1 59840
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output7
timestamp 1
transform 1 0 100188 0 -1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output8
timestamp 1
transform 1 0 100188 0 -1 60928
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp 1
transform -1 0 1748 0 1 62016
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 1
transform -1 0 43608 0 1 101184
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 1
transform -1 0 45540 0 1 101184
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 1
transform 1 0 47748 0 1 101184
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 1
transform 1 0 49680 0 1 101184
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 1
transform -1 0 51336 0 1 101184
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp 1
transform -1 0 53268 0 1 101184
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output16
timestamp 1
transform 1 0 55476 0 1 101184
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output17
timestamp 1
transform 1 0 57408 0 1 101184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_1_Left_577
timestamp 1
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_1_Right_105
timestamp 1
transform -1 0 1932 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_2_Left_106
timestamp 1
transform 1 0 97980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_2_Right_289
timestamp 1
transform -1 0 100832 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_1_Left_395
timestamp 1
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_1_Right_0
timestamp 1
transform -1 0 1932 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_2_Left_107
timestamp 1
transform 1 0 97980 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_2_Right_290
timestamp 1
transform -1 0 100832 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_1_Left_396
timestamp 1
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_1_Right_1
timestamp 1
transform -1 0 1932 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_2_Left_108
timestamp 1
transform 1 0 97980 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_2_Right_291
timestamp 1
transform -1 0 100832 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_1_Left_397
timestamp 1
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_1_Right_2
timestamp 1
transform -1 0 1932 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_2_Left_109
timestamp 1
transform 1 0 97980 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_2_Right_292
timestamp 1
transform -1 0 100832 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_1_Left_398
timestamp 1
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_1_Right_3
timestamp 1
transform -1 0 1932 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_2_Left_110
timestamp 1
transform 1 0 97980 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_2_Right_293
timestamp 1
transform -1 0 100832 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_1_Left_399
timestamp 1
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_1_Right_4
timestamp 1
transform -1 0 1932 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_2_Left_111
timestamp 1
transform 1 0 97980 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_2_Right_294
timestamp 1
transform -1 0 100832 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_1_Left_400
timestamp 1
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_1_Right_5
timestamp 1
transform -1 0 1932 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_2_Left_112
timestamp 1
transform 1 0 97980 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_2_Right_295
timestamp 1
transform -1 0 100832 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_1_Left_401
timestamp 1
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_1_Right_6
timestamp 1
transform -1 0 1932 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_2_Left_113
timestamp 1
transform 1 0 97980 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_2_Right_296
timestamp 1
transform -1 0 100832 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_1_Left_402
timestamp 1
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_1_Right_7
timestamp 1
transform -1 0 1932 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_2_Left_114
timestamp 1
transform 1 0 97980 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_2_Right_297
timestamp 1
transform -1 0 100832 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_1_Left_403
timestamp 1
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_1_Right_8
timestamp 1
transform -1 0 1932 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_2_Left_115
timestamp 1
transform 1 0 97980 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_2_Right_298
timestamp 1
transform -1 0 100832 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_1_Left_404
timestamp 1
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_1_Right_9
timestamp 1
transform -1 0 1932 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_2_Left_116
timestamp 1
transform 1 0 97980 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_2_Right_299
timestamp 1
transform -1 0 100832 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_1_Left_405
timestamp 1
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_1_Right_10
timestamp 1
transform -1 0 1932 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_2_Left_117
timestamp 1
transform 1 0 97980 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_2_Right_300
timestamp 1
transform -1 0 100832 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_1_Left_406
timestamp 1
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_1_Right_11
timestamp 1
transform -1 0 1932 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_2_Left_118
timestamp 1
transform 1 0 97980 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_2_Right_301
timestamp 1
transform -1 0 100832 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_1_Left_407
timestamp 1
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_1_Right_12
timestamp 1
transform -1 0 1932 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_2_Left_119
timestamp 1
transform 1 0 97980 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_2_Right_302
timestamp 1
transform -1 0 100832 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_1_Left_408
timestamp 1
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_1_Right_13
timestamp 1
transform -1 0 1932 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_2_Left_120
timestamp 1
transform 1 0 97980 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_2_Right_303
timestamp 1
transform -1 0 100832 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_1_Left_409
timestamp 1
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_1_Right_14
timestamp 1
transform -1 0 1932 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_2_Left_121
timestamp 1
transform 1 0 97980 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_2_Right_304
timestamp 1
transform -1 0 100832 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_1_Left_410
timestamp 1
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_1_Right_15
timestamp 1
transform -1 0 1932 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_2_Left_122
timestamp 1
transform 1 0 97980 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_2_Right_305
timestamp 1
transform -1 0 100832 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_1_Left_411
timestamp 1
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_1_Right_16
timestamp 1
transform -1 0 1932 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_2_Left_123
timestamp 1
transform 1 0 97980 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_2_Right_306
timestamp 1
transform -1 0 100832 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_1_Left_412
timestamp 1
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_1_Right_17
timestamp 1
transform -1 0 1932 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_2_Left_124
timestamp 1
transform 1 0 97980 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_2_Right_307
timestamp 1
transform -1 0 100832 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_1_Left_413
timestamp 1
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_1_Right_18
timestamp 1
transform -1 0 1932 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_2_Left_125
timestamp 1
transform 1 0 97980 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_2_Right_308
timestamp 1
transform -1 0 100832 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_1_Left_414
timestamp 1
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_1_Right_19
timestamp 1
transform -1 0 1932 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_2_Left_126
timestamp 1
transform 1 0 97980 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_2_Right_309
timestamp 1
transform -1 0 100832 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_1_Left_415
timestamp 1
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_1_Right_20
timestamp 1
transform -1 0 1932 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_2_Left_127
timestamp 1
transform 1 0 97980 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_2_Right_310
timestamp 1
transform -1 0 100832 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_1_Left_416
timestamp 1
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_1_Right_21
timestamp 1
transform -1 0 1932 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_2_Left_128
timestamp 1
transform 1 0 97980 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_2_Right_311
timestamp 1
transform -1 0 100832 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_1_Left_417
timestamp 1
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_1_Right_22
timestamp 1
transform -1 0 1932 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_2_Left_129
timestamp 1
transform 1 0 97980 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_2_Right_312
timestamp 1
transform -1 0 100832 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_1_Left_418
timestamp 1
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_1_Right_23
timestamp 1
transform -1 0 1932 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_2_Left_130
timestamp 1
transform 1 0 97980 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_2_Right_313
timestamp 1
transform -1 0 100832 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_1_Left_419
timestamp 1
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_1_Right_24
timestamp 1
transform -1 0 1932 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_2_Left_131
timestamp 1
transform 1 0 97980 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_2_Right_314
timestamp 1
transform -1 0 100832 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_1_Left_420
timestamp 1
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_1_Right_25
timestamp 1
transform -1 0 1932 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_2_Left_132
timestamp 1
transform 1 0 97980 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_2_Right_315
timestamp 1
transform -1 0 100832 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_1_Left_421
timestamp 1
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_1_Right_26
timestamp 1
transform -1 0 1932 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_2_Left_133
timestamp 1
transform 1 0 97980 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_2_Right_316
timestamp 1
transform -1 0 100832 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_1_Left_422
timestamp 1
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_1_Right_27
timestamp 1
transform -1 0 1932 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_2_Left_134
timestamp 1
transform 1 0 97980 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_2_Right_317
timestamp 1
transform -1 0 100832 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_1_Left_423
timestamp 1
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_1_Right_28
timestamp 1
transform -1 0 1932 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_2_Left_135
timestamp 1
transform 1 0 97980 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_2_Right_318
timestamp 1
transform -1 0 100832 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_1_Left_424
timestamp 1
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_1_Right_29
timestamp 1
transform -1 0 1932 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_2_Left_136
timestamp 1
transform 1 0 97980 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_2_Right_319
timestamp 1
transform -1 0 100832 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_1_Left_425
timestamp 1
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_1_Right_30
timestamp 1
transform -1 0 1932 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_2_Left_137
timestamp 1
transform 1 0 97980 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_2_Right_320
timestamp 1
transform -1 0 100832 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_1_Left_426
timestamp 1
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_1_Right_31
timestamp 1
transform -1 0 1932 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_2_Left_138
timestamp 1
transform 1 0 97980 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_2_Right_321
timestamp 1
transform -1 0 100832 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_1_Left_427
timestamp 1
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_1_Right_32
timestamp 1
transform -1 0 1932 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_2_Left_139
timestamp 1
transform 1 0 97980 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_2_Right_322
timestamp 1
transform -1 0 100832 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_1_Left_428
timestamp 1
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_1_Right_33
timestamp 1
transform -1 0 1932 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_2_Left_140
timestamp 1
transform 1 0 97980 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_2_Right_323
timestamp 1
transform -1 0 100832 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_1_Left_429
timestamp 1
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_1_Right_34
timestamp 1
transform -1 0 1932 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_2_Left_141
timestamp 1
transform 1 0 97980 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_2_Right_324
timestamp 1
transform -1 0 100832 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_1_Left_430
timestamp 1
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_1_Right_35
timestamp 1
transform -1 0 1932 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_2_Left_142
timestamp 1
transform 1 0 97980 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_2_Right_325
timestamp 1
transform -1 0 100832 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_1_Left_431
timestamp 1
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_1_Right_36
timestamp 1
transform -1 0 1932 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_2_Left_143
timestamp 1
transform 1 0 97980 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_2_Right_326
timestamp 1
transform -1 0 100832 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_1_Left_432
timestamp 1
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_1_Right_37
timestamp 1
transform -1 0 1932 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_2_Left_144
timestamp 1
transform 1 0 97980 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_2_Right_327
timestamp 1
transform -1 0 100832 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_1_Left_433
timestamp 1
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_1_Right_38
timestamp 1
transform -1 0 1932 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_2_Left_145
timestamp 1
transform 1 0 97980 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_2_Right_328
timestamp 1
transform -1 0 100832 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_1_Left_434
timestamp 1
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_1_Right_39
timestamp 1
transform -1 0 1932 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_2_Left_146
timestamp 1
transform 1 0 97980 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_2_Right_329
timestamp 1
transform -1 0 100832 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_1_Left_435
timestamp 1
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_1_Right_40
timestamp 1
transform -1 0 1932 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_2_Left_147
timestamp 1
transform 1 0 97980 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_2_Right_330
timestamp 1
transform -1 0 100832 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_1_Left_436
timestamp 1
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_1_Right_41
timestamp 1
transform -1 0 1932 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_2_Left_148
timestamp 1
transform 1 0 97980 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_2_Right_331
timestamp 1
transform -1 0 100832 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_1_Left_437
timestamp 1
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_1_Right_42
timestamp 1
transform -1 0 1932 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_2_Left_149
timestamp 1
transform 1 0 97980 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_2_Right_332
timestamp 1
transform -1 0 100832 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_1_Left_438
timestamp 1
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_1_Right_43
timestamp 1
transform -1 0 1932 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_2_Left_150
timestamp 1
transform 1 0 97980 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_2_Right_333
timestamp 1
transform -1 0 100832 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_1_Left_439
timestamp 1
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_1_Right_44
timestamp 1
transform -1 0 1932 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_2_Left_151
timestamp 1
transform 1 0 97980 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_2_Right_334
timestamp 1
transform -1 0 100832 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_1_Left_440
timestamp 1
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_1_Right_45
timestamp 1
transform -1 0 1932 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_2_Left_152
timestamp 1
transform 1 0 97980 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_2_Right_335
timestamp 1
transform -1 0 100832 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_1_Left_441
timestamp 1
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_1_Right_46
timestamp 1
transform -1 0 1932 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_2_Left_153
timestamp 1
transform 1 0 97980 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_2_Right_336
timestamp 1
transform -1 0 100832 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_1_Left_442
timestamp 1
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_1_Right_47
timestamp 1
transform -1 0 1932 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_2_Left_154
timestamp 1
transform 1 0 97980 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_2_Right_337
timestamp 1
transform -1 0 100832 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_1_Left_443
timestamp 1
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_1_Right_48
timestamp 1
transform -1 0 1932 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_2_Left_155
timestamp 1
transform 1 0 97980 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_2_Right_338
timestamp 1
transform -1 0 100832 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_1_Left_444
timestamp 1
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_1_Right_49
timestamp 1
transform -1 0 1932 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_2_Left_156
timestamp 1
transform 1 0 97980 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_2_Right_339
timestamp 1
transform -1 0 100832 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_1_Left_445
timestamp 1
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_1_Right_50
timestamp 1
transform -1 0 1932 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_2_Left_157
timestamp 1
transform 1 0 97980 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_2_Right_340
timestamp 1
transform -1 0 100832 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_1_Left_446
timestamp 1
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_1_Right_51
timestamp 1
transform -1 0 1932 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_2_Left_158
timestamp 1
transform 1 0 97980 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_2_Right_341
timestamp 1
transform -1 0 100832 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_1_Left_447
timestamp 1
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_1_Right_52
timestamp 1
transform -1 0 1932 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_2_Left_159
timestamp 1
transform 1 0 97980 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_2_Right_342
timestamp 1
transform -1 0 100832 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_1_Left_448
timestamp 1
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_1_Right_53
timestamp 1
transform -1 0 1932 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_2_Left_160
timestamp 1
transform 1 0 97980 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_2_Right_343
timestamp 1
transform -1 0 100832 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_1_Left_449
timestamp 1
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_1_Right_54
timestamp 1
transform -1 0 1932 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_2_Left_161
timestamp 1
transform 1 0 97980 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_2_Right_344
timestamp 1
transform -1 0 100832 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_1_Left_450
timestamp 1
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_1_Right_55
timestamp 1
transform -1 0 1932 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_2_Left_162
timestamp 1
transform 1 0 97980 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_2_Right_345
timestamp 1
transform -1 0 100832 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_1_Left_451
timestamp 1
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_1_Right_56
timestamp 1
transform -1 0 1932 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_2_Left_163
timestamp 1
transform 1 0 97980 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_2_Right_346
timestamp 1
transform -1 0 100832 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_1_Left_452
timestamp 1
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_1_Right_57
timestamp 1
transform -1 0 1932 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_2_Left_164
timestamp 1
transform 1 0 97980 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_2_Right_347
timestamp 1
transform -1 0 100832 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_1_Left_453
timestamp 1
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_1_Right_58
timestamp 1
transform -1 0 1932 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_2_Left_165
timestamp 1
transform 1 0 97980 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_2_Right_348
timestamp 1
transform -1 0 100832 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_1_Left_454
timestamp 1
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_1_Right_59
timestamp 1
transform -1 0 1932 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_2_Left_166
timestamp 1
transform 1 0 97980 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_2_Right_349
timestamp 1
transform -1 0 100832 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_1_Left_455
timestamp 1
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_1_Right_60
timestamp 1
transform -1 0 1932 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_2_Left_167
timestamp 1
transform 1 0 97980 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_2_Right_350
timestamp 1
transform -1 0 100832 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_1_Left_456
timestamp 1
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_1_Right_61
timestamp 1
transform -1 0 1932 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_2_Left_168
timestamp 1
transform 1 0 97980 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_2_Right_351
timestamp 1
transform -1 0 100832 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_1_Left_457
timestamp 1
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_1_Right_62
timestamp 1
transform -1 0 1932 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_2_Left_169
timestamp 1
transform 1 0 97980 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_2_Right_352
timestamp 1
transform -1 0 100832 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_1_Left_458
timestamp 1
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_1_Right_63
timestamp 1
transform -1 0 1932 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_2_Left_170
timestamp 1
transform 1 0 97980 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_2_Right_353
timestamp 1
transform -1 0 100832 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_1_Left_459
timestamp 1
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_1_Right_64
timestamp 1
transform -1 0 1932 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_2_Left_171
timestamp 1
transform 1 0 97980 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_2_Right_354
timestamp 1
transform -1 0 100832 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_1_Left_460
timestamp 1
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_1_Right_65
timestamp 1
transform -1 0 1932 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_2_Left_172
timestamp 1
transform 1 0 97980 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_2_Right_355
timestamp 1
transform -1 0 100832 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_1_Left_461
timestamp 1
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_1_Right_66
timestamp 1
transform -1 0 1932 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_2_Left_173
timestamp 1
transform 1 0 97980 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_2_Right_356
timestamp 1
transform -1 0 100832 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_1_Left_462
timestamp 1
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_1_Right_67
timestamp 1
transform -1 0 1932 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_2_Left_174
timestamp 1
transform 1 0 97980 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_2_Right_357
timestamp 1
transform -1 0 100832 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_1_Left_463
timestamp 1
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_1_Right_68
timestamp 1
transform -1 0 1932 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_2_Left_175
timestamp 1
transform 1 0 97980 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_2_Right_358
timestamp 1
transform -1 0 100832 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_1_Left_464
timestamp 1
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_1_Right_69
timestamp 1
transform -1 0 1932 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_2_Left_176
timestamp 1
transform 1 0 97980 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_2_Right_359
timestamp 1
transform -1 0 100832 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_1_Left_465
timestamp 1
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_1_Right_70
timestamp 1
transform -1 0 1932 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_2_Left_177
timestamp 1
transform 1 0 97980 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_2_Right_360
timestamp 1
transform -1 0 100832 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_1_Left_466
timestamp 1
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_1_Right_71
timestamp 1
transform -1 0 1932 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_2_Left_178
timestamp 1
transform 1 0 97980 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_2_Right_361
timestamp 1
transform -1 0 100832 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_1_Left_467
timestamp 1
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_1_Right_72
timestamp 1
transform -1 0 1932 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_2_Left_179
timestamp 1
transform 1 0 97980 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_2_Right_362
timestamp 1
transform -1 0 100832 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_1_Left_468
timestamp 1
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_1_Right_73
timestamp 1
transform -1 0 1932 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_2_Left_180
timestamp 1
transform 1 0 97980 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_2_Right_363
timestamp 1
transform -1 0 100832 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_1_Left_469
timestamp 1
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_1_Right_74
timestamp 1
transform -1 0 1932 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_2_Left_181
timestamp 1
transform 1 0 97980 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_2_Right_364
timestamp 1
transform -1 0 100832 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_1_Left_470
timestamp 1
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_1_Right_75
timestamp 1
transform -1 0 1932 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_2_Left_182
timestamp 1
transform 1 0 97980 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_2_Right_365
timestamp 1
transform -1 0 100832 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_1_Left_471
timestamp 1
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_1_Right_76
timestamp 1
transform -1 0 1932 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_2_Left_183
timestamp 1
transform 1 0 97980 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_2_Right_366
timestamp 1
transform -1 0 100832 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_1_Left_472
timestamp 1
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_1_Right_77
timestamp 1
transform -1 0 1932 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_2_Left_184
timestamp 1
transform 1 0 97980 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_2_Right_367
timestamp 1
transform -1 0 100832 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_1_Left_473
timestamp 1
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_1_Right_78
timestamp 1
transform -1 0 1932 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_2_Left_185
timestamp 1
transform 1 0 97980 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_2_Right_368
timestamp 1
transform -1 0 100832 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_1_Left_474
timestamp 1
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_1_Right_79
timestamp 1
transform -1 0 1932 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_2_Left_186
timestamp 1
transform 1 0 97980 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_2_Right_369
timestamp 1
transform -1 0 100832 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_1_Left_475
timestamp 1
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_1_Right_80
timestamp 1
transform -1 0 1932 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_2_Left_187
timestamp 1
transform 1 0 97980 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_2_Right_370
timestamp 1
transform -1 0 100832 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_1_Left_476
timestamp 1
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_1_Right_81
timestamp 1
transform -1 0 1932 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_2_Left_188
timestamp 1
transform 1 0 97980 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_2_Right_371
timestamp 1
transform -1 0 100832 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_83_1_Left_477
timestamp 1
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_83_1_Right_82
timestamp 1
transform -1 0 1932 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_83_2_Left_189
timestamp 1
transform 1 0 97980 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_83_2_Right_372
timestamp 1
transform -1 0 100832 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_84_1_Left_478
timestamp 1
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_84_1_Right_83
timestamp 1
transform -1 0 1932 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_84_2_Left_190
timestamp 1
transform 1 0 97980 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_84_2_Right_373
timestamp 1
transform -1 0 100832 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_85_1_Left_479
timestamp 1
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_85_1_Right_84
timestamp 1
transform -1 0 1932 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_85_2_Left_191
timestamp 1
transform 1 0 97980 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_85_2_Right_374
timestamp 1
transform -1 0 100832 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_86_1_Left_480
timestamp 1
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_86_1_Right_85
timestamp 1
transform -1 0 1932 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_86_2_Left_192
timestamp 1
transform 1 0 97980 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_86_2_Right_375
timestamp 1
transform -1 0 100832 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_87_1_Left_481
timestamp 1
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_87_1_Right_86
timestamp 1
transform -1 0 1932 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_87_2_Left_193
timestamp 1
transform 1 0 97980 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_87_2_Right_376
timestamp 1
transform -1 0 100832 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_88_1_Left_482
timestamp 1
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_88_1_Right_87
timestamp 1
transform -1 0 1932 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_88_2_Left_194
timestamp 1
transform 1 0 97980 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_88_2_Right_377
timestamp 1
transform -1 0 100832 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_89_1_Left_483
timestamp 1
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_89_1_Right_88
timestamp 1
transform -1 0 1932 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_89_2_Left_195
timestamp 1
transform 1 0 97980 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_89_2_Right_378
timestamp 1
transform -1 0 100832 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_90_1_Left_484
timestamp 1
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_90_1_Right_89
timestamp 1
transform -1 0 1932 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_90_2_Left_196
timestamp 1
transform 1 0 97980 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_90_2_Right_379
timestamp 1
transform -1 0 100832 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_91_1_Left_485
timestamp 1
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_91_1_Right_90
timestamp 1
transform -1 0 1932 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_91_2_Left_197
timestamp 1
transform 1 0 97980 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_91_2_Right_380
timestamp 1
transform -1 0 100832 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_92_1_Left_486
timestamp 1
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_92_1_Right_91
timestamp 1
transform -1 0 1932 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_92_2_Left_198
timestamp 1
transform 1 0 97980 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_92_2_Right_381
timestamp 1
transform -1 0 100832 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_93_1_Left_487
timestamp 1
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_93_1_Right_92
timestamp 1
transform -1 0 1932 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_93_2_Left_199
timestamp 1
transform 1 0 97980 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_93_2_Right_382
timestamp 1
transform -1 0 100832 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_94_1_Left_488
timestamp 1
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_94_1_Right_93
timestamp 1
transform -1 0 1932 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_94_2_Left_200
timestamp 1
transform 1 0 97980 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_94_2_Right_383
timestamp 1
transform -1 0 100832 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_95_1_Left_489
timestamp 1
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_95_1_Right_94
timestamp 1
transform -1 0 1932 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_95_2_Left_201
timestamp 1
transform 1 0 97980 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_95_2_Right_384
timestamp 1
transform -1 0 100832 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_96_1_Left_490
timestamp 1
transform 1 0 1104 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_96_1_Right_95
timestamp 1
transform -1 0 1932 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_96_2_Left_202
timestamp 1
transform 1 0 97980 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_96_2_Right_385
timestamp 1
transform -1 0 100832 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_97_1_Left_491
timestamp 1
transform 1 0 1104 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_97_1_Right_96
timestamp 1
transform -1 0 1932 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_97_2_Left_203
timestamp 1
transform 1 0 97980 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_97_2_Right_386
timestamp 1
transform -1 0 100832 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_98_1_Left_492
timestamp 1
transform 1 0 1104 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_98_1_Right_97
timestamp 1
transform -1 0 1932 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_98_2_Left_204
timestamp 1
transform 1 0 97980 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_98_2_Right_387
timestamp 1
transform -1 0 100832 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_99_1_Left_493
timestamp 1
transform 1 0 1104 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_99_1_Right_98
timestamp 1
transform -1 0 1932 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_99_2_Left_205
timestamp 1
transform 1 0 97980 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_99_2_Right_388
timestamp 1
transform -1 0 100832 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_100_1_Left_494
timestamp 1
transform 1 0 1104 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_100_1_Right_99
timestamp 1
transform -1 0 1932 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_100_2_Left_206
timestamp 1
transform 1 0 97980 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_100_2_Right_389
timestamp 1
transform -1 0 100832 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_101_1_Left_495
timestamp 1
transform 1 0 1104 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_101_1_Right_100
timestamp 1
transform -1 0 1932 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_101_2_Left_207
timestamp 1
transform 1 0 97980 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_101_2_Right_390
timestamp 1
transform -1 0 100832 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_102_1_Left_496
timestamp 1
transform 1 0 1104 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_102_1_Right_101
timestamp 1
transform -1 0 1932 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_102_2_Left_208
timestamp 1
transform 1 0 97980 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_102_2_Right_391
timestamp 1
transform -1 0 100832 0 1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_103_1_Left_497
timestamp 1
transform 1 0 1104 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_103_1_Right_102
timestamp 1
transform -1 0 1932 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_103_2_Left_209
timestamp 1
transform 1 0 97980 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_103_2_Right_392
timestamp 1
transform -1 0 100832 0 -1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_104_1_Left_498
timestamp 1
transform 1 0 1104 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_104_1_Right_103
timestamp 1
transform -1 0 1932 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_104_2_Left_210
timestamp 1
transform 1 0 97980 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_104_2_Right_393
timestamp 1
transform -1 0 100832 0 1 58752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_105_1_Left_499
timestamp 1
transform 1 0 1104 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_105_1_Right_104
timestamp 1
transform -1 0 1932 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_105_2_Left_211
timestamp 1
transform 1 0 97980 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_105_2_Right_394
timestamp 1
transform -1 0 100832 0 -1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_106_Left_500
timestamp 1
transform 1 0 1104 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_106_Right_212
timestamp 1
transform -1 0 100832 0 1 59840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_107_Left_501
timestamp 1
transform 1 0 1104 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_107_Right_213
timestamp 1
transform -1 0 100832 0 -1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_108_Left_502
timestamp 1
transform 1 0 1104 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_108_Right_214
timestamp 1
transform -1 0 100832 0 1 60928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_109_Left_503
timestamp 1
transform 1 0 1104 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_109_Right_215
timestamp 1
transform -1 0 100832 0 -1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_110_Left_504
timestamp 1
transform 1 0 1104 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_110_Right_216
timestamp 1
transform -1 0 100832 0 1 62016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_111_Left_505
timestamp 1
transform 1 0 1104 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_111_Right_217
timestamp 1
transform -1 0 100832 0 -1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_112_Left_506
timestamp 1
transform 1 0 1104 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_112_Right_218
timestamp 1
transform -1 0 100832 0 1 63104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_113_Left_507
timestamp 1
transform 1 0 1104 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_113_Right_219
timestamp 1
transform -1 0 100832 0 -1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_114_Left_508
timestamp 1
transform 1 0 1104 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_114_Right_220
timestamp 1
transform -1 0 100832 0 1 64192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_115_Left_509
timestamp 1
transform 1 0 1104 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_115_Right_221
timestamp 1
transform -1 0 100832 0 -1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_116_Left_510
timestamp 1
transform 1 0 1104 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_116_Right_222
timestamp 1
transform -1 0 100832 0 1 65280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_117_Left_511
timestamp 1
transform 1 0 1104 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_117_Right_223
timestamp 1
transform -1 0 100832 0 -1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_118_Left_512
timestamp 1
transform 1 0 1104 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_118_Right_224
timestamp 1
transform -1 0 100832 0 1 66368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_119_Left_513
timestamp 1
transform 1 0 1104 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_119_Right_225
timestamp 1
transform -1 0 100832 0 -1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_120_Left_514
timestamp 1
transform 1 0 1104 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_120_Right_226
timestamp 1
transform -1 0 100832 0 1 67456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_121_Left_515
timestamp 1
transform 1 0 1104 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_121_Right_227
timestamp 1
transform -1 0 100832 0 -1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_122_Left_516
timestamp 1
transform 1 0 1104 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_122_Right_228
timestamp 1
transform -1 0 100832 0 1 68544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_123_Left_517
timestamp 1
transform 1 0 1104 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_123_Right_229
timestamp 1
transform -1 0 100832 0 -1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_124_Left_518
timestamp 1
transform 1 0 1104 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_124_Right_230
timestamp 1
transform -1 0 100832 0 1 69632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_125_Left_519
timestamp 1
transform 1 0 1104 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_125_Right_231
timestamp 1
transform -1 0 100832 0 -1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_126_Left_520
timestamp 1
transform 1 0 1104 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_126_Right_232
timestamp 1
transform -1 0 100832 0 1 70720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_127_Left_521
timestamp 1
transform 1 0 1104 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_127_Right_233
timestamp 1
transform -1 0 100832 0 -1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_128_Left_522
timestamp 1
transform 1 0 1104 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_128_Right_234
timestamp 1
transform -1 0 100832 0 1 71808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_129_Left_523
timestamp 1
transform 1 0 1104 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_129_Right_235
timestamp 1
transform -1 0 100832 0 -1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_130_Left_524
timestamp 1
transform 1 0 1104 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_130_Right_236
timestamp 1
transform -1 0 100832 0 1 72896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_131_Left_525
timestamp 1
transform 1 0 1104 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_131_Right_237
timestamp 1
transform -1 0 100832 0 -1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_132_Left_526
timestamp 1
transform 1 0 1104 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_132_Right_238
timestamp 1
transform -1 0 100832 0 1 73984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_133_Left_527
timestamp 1
transform 1 0 1104 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_133_Right_239
timestamp 1
transform -1 0 100832 0 -1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_134_Left_528
timestamp 1
transform 1 0 1104 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_134_Right_240
timestamp 1
transform -1 0 100832 0 1 75072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_135_Left_529
timestamp 1
transform 1 0 1104 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_135_Right_241
timestamp 1
transform -1 0 100832 0 -1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_136_Left_530
timestamp 1
transform 1 0 1104 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_136_Right_242
timestamp 1
transform -1 0 100832 0 1 76160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_137_Left_531
timestamp 1
transform 1 0 1104 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_137_Right_243
timestamp 1
transform -1 0 100832 0 -1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_138_Left_532
timestamp 1
transform 1 0 1104 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_138_Right_244
timestamp 1
transform -1 0 100832 0 1 77248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_139_Left_533
timestamp 1
transform 1 0 1104 0 -1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_139_Right_245
timestamp 1
transform -1 0 100832 0 -1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_140_Left_534
timestamp 1
transform 1 0 1104 0 1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_140_Right_246
timestamp 1
transform -1 0 100832 0 1 78336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_141_Left_535
timestamp 1
transform 1 0 1104 0 -1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_141_Right_247
timestamp 1
transform -1 0 100832 0 -1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_142_Left_536
timestamp 1
transform 1 0 1104 0 1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_142_Right_248
timestamp 1
transform -1 0 100832 0 1 79424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_143_Left_537
timestamp 1
transform 1 0 1104 0 -1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_143_Right_249
timestamp 1
transform -1 0 100832 0 -1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_144_Left_538
timestamp 1
transform 1 0 1104 0 1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_144_Right_250
timestamp 1
transform -1 0 100832 0 1 80512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_145_Left_539
timestamp 1
transform 1 0 1104 0 -1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_145_Right_251
timestamp 1
transform -1 0 100832 0 -1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_146_Left_540
timestamp 1
transform 1 0 1104 0 1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_146_Right_252
timestamp 1
transform -1 0 100832 0 1 81600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_147_Left_541
timestamp 1
transform 1 0 1104 0 -1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_147_Right_253
timestamp 1
transform -1 0 100832 0 -1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_148_Left_542
timestamp 1
transform 1 0 1104 0 1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_148_Right_254
timestamp 1
transform -1 0 100832 0 1 82688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_149_Left_543
timestamp 1
transform 1 0 1104 0 -1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_149_Right_255
timestamp 1
transform -1 0 100832 0 -1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_150_Left_544
timestamp 1
transform 1 0 1104 0 1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_150_Right_256
timestamp 1
transform -1 0 100832 0 1 83776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_151_Left_545
timestamp 1
transform 1 0 1104 0 -1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_151_Right_257
timestamp 1
transform -1 0 100832 0 -1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_152_Left_546
timestamp 1
transform 1 0 1104 0 1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_152_Right_258
timestamp 1
transform -1 0 100832 0 1 84864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_153_Left_547
timestamp 1
transform 1 0 1104 0 -1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_153_Right_259
timestamp 1
transform -1 0 100832 0 -1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_154_Left_548
timestamp 1
transform 1 0 1104 0 1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_154_Right_260
timestamp 1
transform -1 0 100832 0 1 85952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_155_Left_549
timestamp 1
transform 1 0 1104 0 -1 87040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_155_Right_261
timestamp 1
transform -1 0 100832 0 -1 87040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_156_Left_550
timestamp 1
transform 1 0 1104 0 1 87040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_156_Right_262
timestamp 1
transform -1 0 100832 0 1 87040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_157_Left_551
timestamp 1
transform 1 0 1104 0 -1 88128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_157_Right_263
timestamp 1
transform -1 0 100832 0 -1 88128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_158_Left_552
timestamp 1
transform 1 0 1104 0 1 88128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_158_Right_264
timestamp 1
transform -1 0 100832 0 1 88128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_159_Left_553
timestamp 1
transform 1 0 1104 0 -1 89216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_159_Right_265
timestamp 1
transform -1 0 100832 0 -1 89216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_160_Left_554
timestamp 1
transform 1 0 1104 0 1 89216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_160_Right_266
timestamp 1
transform -1 0 100832 0 1 89216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_161_Left_555
timestamp 1
transform 1 0 1104 0 -1 90304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_161_Right_267
timestamp 1
transform -1 0 100832 0 -1 90304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_162_Left_556
timestamp 1
transform 1 0 1104 0 1 90304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_162_Right_268
timestamp 1
transform -1 0 100832 0 1 90304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_163_Left_557
timestamp 1
transform 1 0 1104 0 -1 91392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_163_Right_269
timestamp 1
transform -1 0 100832 0 -1 91392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_164_Left_558
timestamp 1
transform 1 0 1104 0 1 91392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_164_Right_270
timestamp 1
transform -1 0 100832 0 1 91392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_165_Left_559
timestamp 1
transform 1 0 1104 0 -1 92480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_165_Right_271
timestamp 1
transform -1 0 100832 0 -1 92480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_166_Left_560
timestamp 1
transform 1 0 1104 0 1 92480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_166_Right_272
timestamp 1
transform -1 0 100832 0 1 92480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_167_Left_561
timestamp 1
transform 1 0 1104 0 -1 93568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_167_Right_273
timestamp 1
transform -1 0 100832 0 -1 93568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_168_Left_562
timestamp 1
transform 1 0 1104 0 1 93568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_168_Right_274
timestamp 1
transform -1 0 100832 0 1 93568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_169_Left_563
timestamp 1
transform 1 0 1104 0 -1 94656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_169_Right_275
timestamp 1
transform -1 0 100832 0 -1 94656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_170_Left_564
timestamp 1
transform 1 0 1104 0 1 94656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_170_Right_276
timestamp 1
transform -1 0 100832 0 1 94656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_171_Left_565
timestamp 1
transform 1 0 1104 0 -1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_171_Right_277
timestamp 1
transform -1 0 100832 0 -1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_172_Left_566
timestamp 1
transform 1 0 1104 0 1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_172_Right_278
timestamp 1
transform -1 0 100832 0 1 95744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_173_Left_567
timestamp 1
transform 1 0 1104 0 -1 96832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_173_Right_279
timestamp 1
transform -1 0 100832 0 -1 96832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_174_Left_568
timestamp 1
transform 1 0 1104 0 1 96832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_174_Right_280
timestamp 1
transform -1 0 100832 0 1 96832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_175_Left_569
timestamp 1
transform 1 0 1104 0 -1 97920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_175_Right_281
timestamp 1
transform -1 0 100832 0 -1 97920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_176_Left_570
timestamp 1
transform 1 0 1104 0 1 97920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_176_Right_282
timestamp 1
transform -1 0 100832 0 1 97920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_177_Left_571
timestamp 1
transform 1 0 1104 0 -1 99008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_177_Right_283
timestamp 1
transform -1 0 100832 0 -1 99008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_178_Left_572
timestamp 1
transform 1 0 1104 0 1 99008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_178_Right_284
timestamp 1
transform -1 0 100832 0 1 99008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_179_Left_573
timestamp 1
transform 1 0 1104 0 -1 100096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_179_Right_285
timestamp 1
transform -1 0 100832 0 -1 100096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_180_Left_574
timestamp 1
transform 1 0 1104 0 1 100096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_180_Right_286
timestamp 1
transform -1 0 100832 0 1 100096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_181_Left_575
timestamp 1
transform 1 0 1104 0 -1 101184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_181_Right_287
timestamp 1
transform -1 0 100832 0 -1 101184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_182_Left_576
timestamp 1
transform 1 0 1104 0 1 101184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_182_Right_288
timestamp 1
transform -1 0 100832 0 1 101184
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_578
timestamp 1
transform 1 0 3680 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_579
timestamp 1
transform 1 0 6256 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_580
timestamp 1
transform 1 0 8832 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_581
timestamp 1
transform 1 0 11408 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_582
timestamp 1
transform 1 0 13984 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_583
timestamp 1
transform 1 0 16560 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_584
timestamp 1
transform 1 0 19136 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_585
timestamp 1
transform 1 0 21712 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_586
timestamp 1
transform 1 0 24288 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_587
timestamp 1
transform 1 0 26864 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_588
timestamp 1
transform 1 0 29440 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_589
timestamp 1
transform 1 0 32016 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_590
timestamp 1
transform 1 0 34592 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_591
timestamp 1
transform 1 0 37168 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_592
timestamp 1
transform 1 0 39744 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_593
timestamp 1
transform 1 0 42320 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_594
timestamp 1
transform 1 0 44896 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_595
timestamp 1
transform 1 0 47472 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_596
timestamp 1
transform 1 0 50048 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_597
timestamp 1
transform 1 0 52624 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_598
timestamp 1
transform 1 0 55200 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_599
timestamp 1
transform 1 0 57776 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_600
timestamp 1
transform 1 0 60352 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_601
timestamp 1
transform 1 0 62928 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_602
timestamp 1
transform 1 0 65504 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_603
timestamp 1
transform 1 0 68080 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_604
timestamp 1
transform 1 0 70656 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_605
timestamp 1
transform 1 0 73232 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_606
timestamp 1
transform 1 0 75808 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_607
timestamp 1
transform 1 0 78384 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_608
timestamp 1
transform 1 0 80960 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_609
timestamp 1
transform 1 0 83536 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_610
timestamp 1
transform 1 0 86112 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_611
timestamp 1
transform 1 0 88688 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_612
timestamp 1
transform 1 0 91264 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_613
timestamp 1
transform 1 0 93840 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_614
timestamp 1
transform 1 0 96416 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_615
timestamp 1
transform 1 0 98992 0 1 59840
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_107_616
timestamp 1
transform 1 0 6256 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_107_617
timestamp 1
transform 1 0 11408 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_107_618
timestamp 1
transform 1 0 16560 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_107_619
timestamp 1
transform 1 0 21712 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_107_620
timestamp 1
transform 1 0 26864 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_107_621
timestamp 1
transform 1 0 32016 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_107_622
timestamp 1
transform 1 0 37168 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_107_623
timestamp 1
transform 1 0 42320 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_107_624
timestamp 1
transform 1 0 47472 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_107_625
timestamp 1
transform 1 0 52624 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_107_626
timestamp 1
transform 1 0 57776 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_107_627
timestamp 1
transform 1 0 62928 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_107_628
timestamp 1
transform 1 0 68080 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_107_629
timestamp 1
transform 1 0 73232 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_107_630
timestamp 1
transform 1 0 78384 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_107_631
timestamp 1
transform 1 0 83536 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_107_632
timestamp 1
transform 1 0 88688 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_107_633
timestamp 1
transform 1 0 93840 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_107_634
timestamp 1
transform 1 0 98992 0 -1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_635
timestamp 1
transform 1 0 3680 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_636
timestamp 1
transform 1 0 8832 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_637
timestamp 1
transform 1 0 13984 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_638
timestamp 1
transform 1 0 19136 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_639
timestamp 1
transform 1 0 24288 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_640
timestamp 1
transform 1 0 29440 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_641
timestamp 1
transform 1 0 34592 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_642
timestamp 1
transform 1 0 39744 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_643
timestamp 1
transform 1 0 44896 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_644
timestamp 1
transform 1 0 50048 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_645
timestamp 1
transform 1 0 55200 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_646
timestamp 1
transform 1 0 60352 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_647
timestamp 1
transform 1 0 65504 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_648
timestamp 1
transform 1 0 70656 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_649
timestamp 1
transform 1 0 75808 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_650
timestamp 1
transform 1 0 80960 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_651
timestamp 1
transform 1 0 86112 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_652
timestamp 1
transform 1 0 91264 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_653
timestamp 1
transform 1 0 96416 0 1 60928
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_109_654
timestamp 1
transform 1 0 6256 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_109_655
timestamp 1
transform 1 0 11408 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_109_656
timestamp 1
transform 1 0 16560 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_109_657
timestamp 1
transform 1 0 21712 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_109_658
timestamp 1
transform 1 0 26864 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_109_659
timestamp 1
transform 1 0 32016 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_109_660
timestamp 1
transform 1 0 37168 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_109_661
timestamp 1
transform 1 0 42320 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_109_662
timestamp 1
transform 1 0 47472 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_109_663
timestamp 1
transform 1 0 52624 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_109_664
timestamp 1
transform 1 0 57776 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_109_665
timestamp 1
transform 1 0 62928 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_109_666
timestamp 1
transform 1 0 68080 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_109_667
timestamp 1
transform 1 0 73232 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_109_668
timestamp 1
transform 1 0 78384 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_109_669
timestamp 1
transform 1 0 83536 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_109_670
timestamp 1
transform 1 0 88688 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_109_671
timestamp 1
transform 1 0 93840 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_109_672
timestamp 1
transform 1 0 98992 0 -1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_673
timestamp 1
transform 1 0 3680 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_674
timestamp 1
transform 1 0 8832 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_675
timestamp 1
transform 1 0 13984 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_676
timestamp 1
transform 1 0 19136 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_677
timestamp 1
transform 1 0 24288 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_678
timestamp 1
transform 1 0 29440 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_679
timestamp 1
transform 1 0 34592 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_680
timestamp 1
transform 1 0 39744 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_681
timestamp 1
transform 1 0 44896 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_682
timestamp 1
transform 1 0 50048 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_683
timestamp 1
transform 1 0 55200 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_684
timestamp 1
transform 1 0 60352 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_685
timestamp 1
transform 1 0 65504 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_686
timestamp 1
transform 1 0 70656 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_687
timestamp 1
transform 1 0 75808 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_688
timestamp 1
transform 1 0 80960 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_689
timestamp 1
transform 1 0 86112 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_690
timestamp 1
transform 1 0 91264 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_691
timestamp 1
transform 1 0 96416 0 1 62016
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_111_692
timestamp 1
transform 1 0 6256 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_111_693
timestamp 1
transform 1 0 11408 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_111_694
timestamp 1
transform 1 0 16560 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_111_695
timestamp 1
transform 1 0 21712 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_111_696
timestamp 1
transform 1 0 26864 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_111_697
timestamp 1
transform 1 0 32016 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_111_698
timestamp 1
transform 1 0 37168 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_111_699
timestamp 1
transform 1 0 42320 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_111_700
timestamp 1
transform 1 0 47472 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_111_701
timestamp 1
transform 1 0 52624 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_111_702
timestamp 1
transform 1 0 57776 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_111_703
timestamp 1
transform 1 0 62928 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_111_704
timestamp 1
transform 1 0 68080 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_111_705
timestamp 1
transform 1 0 73232 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_111_706
timestamp 1
transform 1 0 78384 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_111_707
timestamp 1
transform 1 0 83536 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_111_708
timestamp 1
transform 1 0 88688 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_111_709
timestamp 1
transform 1 0 93840 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_111_710
timestamp 1
transform 1 0 98992 0 -1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_711
timestamp 1
transform 1 0 3680 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_712
timestamp 1
transform 1 0 8832 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_713
timestamp 1
transform 1 0 13984 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_714
timestamp 1
transform 1 0 19136 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_715
timestamp 1
transform 1 0 24288 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_716
timestamp 1
transform 1 0 29440 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_717
timestamp 1
transform 1 0 34592 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_718
timestamp 1
transform 1 0 39744 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_719
timestamp 1
transform 1 0 44896 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_720
timestamp 1
transform 1 0 50048 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_721
timestamp 1
transform 1 0 55200 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_722
timestamp 1
transform 1 0 60352 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_723
timestamp 1
transform 1 0 65504 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_724
timestamp 1
transform 1 0 70656 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_725
timestamp 1
transform 1 0 75808 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_726
timestamp 1
transform 1 0 80960 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_727
timestamp 1
transform 1 0 86112 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_728
timestamp 1
transform 1 0 91264 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_729
timestamp 1
transform 1 0 96416 0 1 63104
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_113_730
timestamp 1
transform 1 0 6256 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_113_731
timestamp 1
transform 1 0 11408 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_113_732
timestamp 1
transform 1 0 16560 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_113_733
timestamp 1
transform 1 0 21712 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_113_734
timestamp 1
transform 1 0 26864 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_113_735
timestamp 1
transform 1 0 32016 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_113_736
timestamp 1
transform 1 0 37168 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_113_737
timestamp 1
transform 1 0 42320 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_113_738
timestamp 1
transform 1 0 47472 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_113_739
timestamp 1
transform 1 0 52624 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_113_740
timestamp 1
transform 1 0 57776 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_113_741
timestamp 1
transform 1 0 62928 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_113_742
timestamp 1
transform 1 0 68080 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_113_743
timestamp 1
transform 1 0 73232 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_113_744
timestamp 1
transform 1 0 78384 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_113_745
timestamp 1
transform 1 0 83536 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_113_746
timestamp 1
transform 1 0 88688 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_113_747
timestamp 1
transform 1 0 93840 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_113_748
timestamp 1
transform 1 0 98992 0 -1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_749
timestamp 1
transform 1 0 3680 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_750
timestamp 1
transform 1 0 8832 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_751
timestamp 1
transform 1 0 13984 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_752
timestamp 1
transform 1 0 19136 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_753
timestamp 1
transform 1 0 24288 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_754
timestamp 1
transform 1 0 29440 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_755
timestamp 1
transform 1 0 34592 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_756
timestamp 1
transform 1 0 39744 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_757
timestamp 1
transform 1 0 44896 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_758
timestamp 1
transform 1 0 50048 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_759
timestamp 1
transform 1 0 55200 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_760
timestamp 1
transform 1 0 60352 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_761
timestamp 1
transform 1 0 65504 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_762
timestamp 1
transform 1 0 70656 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_763
timestamp 1
transform 1 0 75808 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_764
timestamp 1
transform 1 0 80960 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_765
timestamp 1
transform 1 0 86112 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_766
timestamp 1
transform 1 0 91264 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_767
timestamp 1
transform 1 0 96416 0 1 64192
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_115_768
timestamp 1
transform 1 0 6256 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_115_769
timestamp 1
transform 1 0 11408 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_115_770
timestamp 1
transform 1 0 16560 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_115_771
timestamp 1
transform 1 0 21712 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_115_772
timestamp 1
transform 1 0 26864 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_115_773
timestamp 1
transform 1 0 32016 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_115_774
timestamp 1
transform 1 0 37168 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_115_775
timestamp 1
transform 1 0 42320 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_115_776
timestamp 1
transform 1 0 47472 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_115_777
timestamp 1
transform 1 0 52624 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_115_778
timestamp 1
transform 1 0 57776 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_115_779
timestamp 1
transform 1 0 62928 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_115_780
timestamp 1
transform 1 0 68080 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_115_781
timestamp 1
transform 1 0 73232 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_115_782
timestamp 1
transform 1 0 78384 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_115_783
timestamp 1
transform 1 0 83536 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_115_784
timestamp 1
transform 1 0 88688 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_115_785
timestamp 1
transform 1 0 93840 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_115_786
timestamp 1
transform 1 0 98992 0 -1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_787
timestamp 1
transform 1 0 3680 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_788
timestamp 1
transform 1 0 8832 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_789
timestamp 1
transform 1 0 13984 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_790
timestamp 1
transform 1 0 19136 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_791
timestamp 1
transform 1 0 24288 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_792
timestamp 1
transform 1 0 29440 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_793
timestamp 1
transform 1 0 34592 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_794
timestamp 1
transform 1 0 39744 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_795
timestamp 1
transform 1 0 44896 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_796
timestamp 1
transform 1 0 50048 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_797
timestamp 1
transform 1 0 55200 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_798
timestamp 1
transform 1 0 60352 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_799
timestamp 1
transform 1 0 65504 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_800
timestamp 1
transform 1 0 70656 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_801
timestamp 1
transform 1 0 75808 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_802
timestamp 1
transform 1 0 80960 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_803
timestamp 1
transform 1 0 86112 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_804
timestamp 1
transform 1 0 91264 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_805
timestamp 1
transform 1 0 96416 0 1 65280
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_806
timestamp 1
transform 1 0 6256 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_807
timestamp 1
transform 1 0 11408 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_808
timestamp 1
transform 1 0 16560 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_809
timestamp 1
transform 1 0 21712 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_810
timestamp 1
transform 1 0 26864 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_811
timestamp 1
transform 1 0 32016 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_812
timestamp 1
transform 1 0 37168 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_813
timestamp 1
transform 1 0 42320 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_814
timestamp 1
transform 1 0 47472 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_815
timestamp 1
transform 1 0 52624 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_816
timestamp 1
transform 1 0 57776 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_817
timestamp 1
transform 1 0 62928 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_818
timestamp 1
transform 1 0 68080 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_819
timestamp 1
transform 1 0 73232 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_820
timestamp 1
transform 1 0 78384 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_821
timestamp 1
transform 1 0 83536 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_822
timestamp 1
transform 1 0 88688 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_823
timestamp 1
transform 1 0 93840 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_117_824
timestamp 1
transform 1 0 98992 0 -1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_825
timestamp 1
transform 1 0 3680 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_826
timestamp 1
transform 1 0 8832 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_827
timestamp 1
transform 1 0 13984 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_828
timestamp 1
transform 1 0 19136 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_829
timestamp 1
transform 1 0 24288 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_830
timestamp 1
transform 1 0 29440 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_831
timestamp 1
transform 1 0 34592 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_832
timestamp 1
transform 1 0 39744 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_833
timestamp 1
transform 1 0 44896 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_834
timestamp 1
transform 1 0 50048 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_835
timestamp 1
transform 1 0 55200 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_836
timestamp 1
transform 1 0 60352 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_837
timestamp 1
transform 1 0 65504 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_838
timestamp 1
transform 1 0 70656 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_839
timestamp 1
transform 1 0 75808 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_840
timestamp 1
transform 1 0 80960 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_841
timestamp 1
transform 1 0 86112 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_842
timestamp 1
transform 1 0 91264 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_843
timestamp 1
transform 1 0 96416 0 1 66368
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_844
timestamp 1
transform 1 0 6256 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_845
timestamp 1
transform 1 0 11408 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_846
timestamp 1
transform 1 0 16560 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_847
timestamp 1
transform 1 0 21712 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_848
timestamp 1
transform 1 0 26864 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_849
timestamp 1
transform 1 0 32016 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_850
timestamp 1
transform 1 0 37168 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_851
timestamp 1
transform 1 0 42320 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_852
timestamp 1
transform 1 0 47472 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_853
timestamp 1
transform 1 0 52624 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_854
timestamp 1
transform 1 0 57776 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_855
timestamp 1
transform 1 0 62928 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_856
timestamp 1
transform 1 0 68080 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_857
timestamp 1
transform 1 0 73232 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_858
timestamp 1
transform 1 0 78384 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_859
timestamp 1
transform 1 0 83536 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_860
timestamp 1
transform 1 0 88688 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_861
timestamp 1
transform 1 0 93840 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_119_862
timestamp 1
transform 1 0 98992 0 -1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_863
timestamp 1
transform 1 0 3680 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_864
timestamp 1
transform 1 0 8832 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_865
timestamp 1
transform 1 0 13984 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_866
timestamp 1
transform 1 0 19136 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_867
timestamp 1
transform 1 0 24288 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_868
timestamp 1
transform 1 0 29440 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_869
timestamp 1
transform 1 0 34592 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_870
timestamp 1
transform 1 0 39744 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_871
timestamp 1
transform 1 0 44896 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_872
timestamp 1
transform 1 0 50048 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_873
timestamp 1
transform 1 0 55200 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_874
timestamp 1
transform 1 0 60352 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_875
timestamp 1
transform 1 0 65504 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_876
timestamp 1
transform 1 0 70656 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_877
timestamp 1
transform 1 0 75808 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_878
timestamp 1
transform 1 0 80960 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_879
timestamp 1
transform 1 0 86112 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_880
timestamp 1
transform 1 0 91264 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_881
timestamp 1
transform 1 0 96416 0 1 67456
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_882
timestamp 1
transform 1 0 6256 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_883
timestamp 1
transform 1 0 11408 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_884
timestamp 1
transform 1 0 16560 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_885
timestamp 1
transform 1 0 21712 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_886
timestamp 1
transform 1 0 26864 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_887
timestamp 1
transform 1 0 32016 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_888
timestamp 1
transform 1 0 37168 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_889
timestamp 1
transform 1 0 42320 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_890
timestamp 1
transform 1 0 47472 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_891
timestamp 1
transform 1 0 52624 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_892
timestamp 1
transform 1 0 57776 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_893
timestamp 1
transform 1 0 62928 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_894
timestamp 1
transform 1 0 68080 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_895
timestamp 1
transform 1 0 73232 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_896
timestamp 1
transform 1 0 78384 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_897
timestamp 1
transform 1 0 83536 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_898
timestamp 1
transform 1 0 88688 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_899
timestamp 1
transform 1 0 93840 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_121_900
timestamp 1
transform 1 0 98992 0 -1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_901
timestamp 1
transform 1 0 3680 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_902
timestamp 1
transform 1 0 8832 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_903
timestamp 1
transform 1 0 13984 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_904
timestamp 1
transform 1 0 19136 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_905
timestamp 1
transform 1 0 24288 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_906
timestamp 1
transform 1 0 29440 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_907
timestamp 1
transform 1 0 34592 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_908
timestamp 1
transform 1 0 39744 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_909
timestamp 1
transform 1 0 44896 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_910
timestamp 1
transform 1 0 50048 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_911
timestamp 1
transform 1 0 55200 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_912
timestamp 1
transform 1 0 60352 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_913
timestamp 1
transform 1 0 65504 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_914
timestamp 1
transform 1 0 70656 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_915
timestamp 1
transform 1 0 75808 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_916
timestamp 1
transform 1 0 80960 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_917
timestamp 1
transform 1 0 86112 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_918
timestamp 1
transform 1 0 91264 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_919
timestamp 1
transform 1 0 96416 0 1 68544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_920
timestamp 1
transform 1 0 6256 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_921
timestamp 1
transform 1 0 11408 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_922
timestamp 1
transform 1 0 16560 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_923
timestamp 1
transform 1 0 21712 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_924
timestamp 1
transform 1 0 26864 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_925
timestamp 1
transform 1 0 32016 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_926
timestamp 1
transform 1 0 37168 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_927
timestamp 1
transform 1 0 42320 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_928
timestamp 1
transform 1 0 47472 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_929
timestamp 1
transform 1 0 52624 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_930
timestamp 1
transform 1 0 57776 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_931
timestamp 1
transform 1 0 62928 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_932
timestamp 1
transform 1 0 68080 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_933
timestamp 1
transform 1 0 73232 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_934
timestamp 1
transform 1 0 78384 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_935
timestamp 1
transform 1 0 83536 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_936
timestamp 1
transform 1 0 88688 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_937
timestamp 1
transform 1 0 93840 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_123_938
timestamp 1
transform 1 0 98992 0 -1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_939
timestamp 1
transform 1 0 3680 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_940
timestamp 1
transform 1 0 8832 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_941
timestamp 1
transform 1 0 13984 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_942
timestamp 1
transform 1 0 19136 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_943
timestamp 1
transform 1 0 24288 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_944
timestamp 1
transform 1 0 29440 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_945
timestamp 1
transform 1 0 34592 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_946
timestamp 1
transform 1 0 39744 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_947
timestamp 1
transform 1 0 44896 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_948
timestamp 1
transform 1 0 50048 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_949
timestamp 1
transform 1 0 55200 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_950
timestamp 1
transform 1 0 60352 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_951
timestamp 1
transform 1 0 65504 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_952
timestamp 1
transform 1 0 70656 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_953
timestamp 1
transform 1 0 75808 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_954
timestamp 1
transform 1 0 80960 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_955
timestamp 1
transform 1 0 86112 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_956
timestamp 1
transform 1 0 91264 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_957
timestamp 1
transform 1 0 96416 0 1 69632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_958
timestamp 1
transform 1 0 6256 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_959
timestamp 1
transform 1 0 11408 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_960
timestamp 1
transform 1 0 16560 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_961
timestamp 1
transform 1 0 21712 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_962
timestamp 1
transform 1 0 26864 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_963
timestamp 1
transform 1 0 32016 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_964
timestamp 1
transform 1 0 37168 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_965
timestamp 1
transform 1 0 42320 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_966
timestamp 1
transform 1 0 47472 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_967
timestamp 1
transform 1 0 52624 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_968
timestamp 1
transform 1 0 57776 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_969
timestamp 1
transform 1 0 62928 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_970
timestamp 1
transform 1 0 68080 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_971
timestamp 1
transform 1 0 73232 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_972
timestamp 1
transform 1 0 78384 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_973
timestamp 1
transform 1 0 83536 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_974
timestamp 1
transform 1 0 88688 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_975
timestamp 1
transform 1 0 93840 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_125_976
timestamp 1
transform 1 0 98992 0 -1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_977
timestamp 1
transform 1 0 3680 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_978
timestamp 1
transform 1 0 8832 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_979
timestamp 1
transform 1 0 13984 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_980
timestamp 1
transform 1 0 19136 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_981
timestamp 1
transform 1 0 24288 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_982
timestamp 1
transform 1 0 29440 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_983
timestamp 1
transform 1 0 34592 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_984
timestamp 1
transform 1 0 39744 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_985
timestamp 1
transform 1 0 44896 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_986
timestamp 1
transform 1 0 50048 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_987
timestamp 1
transform 1 0 55200 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_988
timestamp 1
transform 1 0 60352 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_989
timestamp 1
transform 1 0 65504 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_990
timestamp 1
transform 1 0 70656 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_991
timestamp 1
transform 1 0 75808 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_992
timestamp 1
transform 1 0 80960 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_993
timestamp 1
transform 1 0 86112 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_994
timestamp 1
transform 1 0 91264 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_995
timestamp 1
transform 1 0 96416 0 1 70720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_996
timestamp 1
transform 1 0 6256 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_997
timestamp 1
transform 1 0 11408 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_998
timestamp 1
transform 1 0 16560 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_999
timestamp 1
transform 1 0 21712 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1000
timestamp 1
transform 1 0 26864 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1001
timestamp 1
transform 1 0 32016 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1002
timestamp 1
transform 1 0 37168 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1003
timestamp 1
transform 1 0 42320 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1004
timestamp 1
transform 1 0 47472 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1005
timestamp 1
transform 1 0 52624 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1006
timestamp 1
transform 1 0 57776 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1007
timestamp 1
transform 1 0 62928 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1008
timestamp 1
transform 1 0 68080 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1009
timestamp 1
transform 1 0 73232 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1010
timestamp 1
transform 1 0 78384 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1011
timestamp 1
transform 1 0 83536 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1012
timestamp 1
transform 1 0 88688 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1013
timestamp 1
transform 1 0 93840 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_127_1014
timestamp 1
transform 1 0 98992 0 -1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_1015
timestamp 1
transform 1 0 3680 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_1016
timestamp 1
transform 1 0 8832 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_1017
timestamp 1
transform 1 0 13984 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_1018
timestamp 1
transform 1 0 19136 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_1019
timestamp 1
transform 1 0 24288 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_1020
timestamp 1
transform 1 0 29440 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_1021
timestamp 1
transform 1 0 34592 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_1022
timestamp 1
transform 1 0 39744 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_1023
timestamp 1
transform 1 0 44896 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_1024
timestamp 1
transform 1 0 50048 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_1025
timestamp 1
transform 1 0 55200 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_1026
timestamp 1
transform 1 0 60352 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_1027
timestamp 1
transform 1 0 65504 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_1028
timestamp 1
transform 1 0 70656 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_1029
timestamp 1
transform 1 0 75808 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_1030
timestamp 1
transform 1 0 80960 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_1031
timestamp 1
transform 1 0 86112 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_1032
timestamp 1
transform 1 0 91264 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_1033
timestamp 1
transform 1 0 96416 0 1 71808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_1034
timestamp 1
transform 1 0 6256 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_1035
timestamp 1
transform 1 0 11408 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_1036
timestamp 1
transform 1 0 16560 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_1037
timestamp 1
transform 1 0 21712 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_1038
timestamp 1
transform 1 0 26864 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_1039
timestamp 1
transform 1 0 32016 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_1040
timestamp 1
transform 1 0 37168 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_1041
timestamp 1
transform 1 0 42320 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_1042
timestamp 1
transform 1 0 47472 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_1043
timestamp 1
transform 1 0 52624 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_1044
timestamp 1
transform 1 0 57776 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_1045
timestamp 1
transform 1 0 62928 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_1046
timestamp 1
transform 1 0 68080 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_1047
timestamp 1
transform 1 0 73232 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_1048
timestamp 1
transform 1 0 78384 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_1049
timestamp 1
transform 1 0 83536 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_1050
timestamp 1
transform 1 0 88688 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_1051
timestamp 1
transform 1 0 93840 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_129_1052
timestamp 1
transform 1 0 98992 0 -1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_1053
timestamp 1
transform 1 0 3680 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_1054
timestamp 1
transform 1 0 8832 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_1055
timestamp 1
transform 1 0 13984 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_1056
timestamp 1
transform 1 0 19136 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_1057
timestamp 1
transform 1 0 24288 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_1058
timestamp 1
transform 1 0 29440 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_1059
timestamp 1
transform 1 0 34592 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_1060
timestamp 1
transform 1 0 39744 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_1061
timestamp 1
transform 1 0 44896 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_1062
timestamp 1
transform 1 0 50048 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_1063
timestamp 1
transform 1 0 55200 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_1064
timestamp 1
transform 1 0 60352 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_1065
timestamp 1
transform 1 0 65504 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_1066
timestamp 1
transform 1 0 70656 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_1067
timestamp 1
transform 1 0 75808 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_1068
timestamp 1
transform 1 0 80960 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_1069
timestamp 1
transform 1 0 86112 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_1070
timestamp 1
transform 1 0 91264 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_1071
timestamp 1
transform 1 0 96416 0 1 72896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_1072
timestamp 1
transform 1 0 6256 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_1073
timestamp 1
transform 1 0 11408 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_1074
timestamp 1
transform 1 0 16560 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_1075
timestamp 1
transform 1 0 21712 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_1076
timestamp 1
transform 1 0 26864 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_1077
timestamp 1
transform 1 0 32016 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_1078
timestamp 1
transform 1 0 37168 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_1079
timestamp 1
transform 1 0 42320 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_1080
timestamp 1
transform 1 0 47472 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_1081
timestamp 1
transform 1 0 52624 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_1082
timestamp 1
transform 1 0 57776 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_1083
timestamp 1
transform 1 0 62928 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_1084
timestamp 1
transform 1 0 68080 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_1085
timestamp 1
transform 1 0 73232 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_1086
timestamp 1
transform 1 0 78384 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_1087
timestamp 1
transform 1 0 83536 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_1088
timestamp 1
transform 1 0 88688 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_1089
timestamp 1
transform 1 0 93840 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_131_1090
timestamp 1
transform 1 0 98992 0 -1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_1091
timestamp 1
transform 1 0 3680 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_1092
timestamp 1
transform 1 0 8832 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_1093
timestamp 1
transform 1 0 13984 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_1094
timestamp 1
transform 1 0 19136 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_1095
timestamp 1
transform 1 0 24288 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_1096
timestamp 1
transform 1 0 29440 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_1097
timestamp 1
transform 1 0 34592 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_1098
timestamp 1
transform 1 0 39744 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_1099
timestamp 1
transform 1 0 44896 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_1100
timestamp 1
transform 1 0 50048 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_1101
timestamp 1
transform 1 0 55200 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_1102
timestamp 1
transform 1 0 60352 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_1103
timestamp 1
transform 1 0 65504 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_1104
timestamp 1
transform 1 0 70656 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_1105
timestamp 1
transform 1 0 75808 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_1106
timestamp 1
transform 1 0 80960 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_1107
timestamp 1
transform 1 0 86112 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_1108
timestamp 1
transform 1 0 91264 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_1109
timestamp 1
transform 1 0 96416 0 1 73984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_1110
timestamp 1
transform 1 0 6256 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_1111
timestamp 1
transform 1 0 11408 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_1112
timestamp 1
transform 1 0 16560 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_1113
timestamp 1
transform 1 0 21712 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_1114
timestamp 1
transform 1 0 26864 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_1115
timestamp 1
transform 1 0 32016 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_1116
timestamp 1
transform 1 0 37168 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_1117
timestamp 1
transform 1 0 42320 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_1118
timestamp 1
transform 1 0 47472 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_1119
timestamp 1
transform 1 0 52624 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_1120
timestamp 1
transform 1 0 57776 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_1121
timestamp 1
transform 1 0 62928 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_1122
timestamp 1
transform 1 0 68080 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_1123
timestamp 1
transform 1 0 73232 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_1124
timestamp 1
transform 1 0 78384 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_1125
timestamp 1
transform 1 0 83536 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_1126
timestamp 1
transform 1 0 88688 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_1127
timestamp 1
transform 1 0 93840 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_133_1128
timestamp 1
transform 1 0 98992 0 -1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_1129
timestamp 1
transform 1 0 3680 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_1130
timestamp 1
transform 1 0 8832 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_1131
timestamp 1
transform 1 0 13984 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_1132
timestamp 1
transform 1 0 19136 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_1133
timestamp 1
transform 1 0 24288 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_1134
timestamp 1
transform 1 0 29440 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_1135
timestamp 1
transform 1 0 34592 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_1136
timestamp 1
transform 1 0 39744 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_1137
timestamp 1
transform 1 0 44896 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_1138
timestamp 1
transform 1 0 50048 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_1139
timestamp 1
transform 1 0 55200 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_1140
timestamp 1
transform 1 0 60352 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_1141
timestamp 1
transform 1 0 65504 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_1142
timestamp 1
transform 1 0 70656 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_1143
timestamp 1
transform 1 0 75808 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_1144
timestamp 1
transform 1 0 80960 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_1145
timestamp 1
transform 1 0 86112 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_1146
timestamp 1
transform 1 0 91264 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_1147
timestamp 1
transform 1 0 96416 0 1 75072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_1148
timestamp 1
transform 1 0 6256 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_1149
timestamp 1
transform 1 0 11408 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_1150
timestamp 1
transform 1 0 16560 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_1151
timestamp 1
transform 1 0 21712 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_1152
timestamp 1
transform 1 0 26864 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_1153
timestamp 1
transform 1 0 32016 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_1154
timestamp 1
transform 1 0 37168 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_1155
timestamp 1
transform 1 0 42320 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_1156
timestamp 1
transform 1 0 47472 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_1157
timestamp 1
transform 1 0 52624 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_1158
timestamp 1
transform 1 0 57776 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_1159
timestamp 1
transform 1 0 62928 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_1160
timestamp 1
transform 1 0 68080 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_1161
timestamp 1
transform 1 0 73232 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_1162
timestamp 1
transform 1 0 78384 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_1163
timestamp 1
transform 1 0 83536 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_1164
timestamp 1
transform 1 0 88688 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_1165
timestamp 1
transform 1 0 93840 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_135_1166
timestamp 1
transform 1 0 98992 0 -1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_1167
timestamp 1
transform 1 0 3680 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_1168
timestamp 1
transform 1 0 8832 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_1169
timestamp 1
transform 1 0 13984 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_1170
timestamp 1
transform 1 0 19136 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_1171
timestamp 1
transform 1 0 24288 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_1172
timestamp 1
transform 1 0 29440 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_1173
timestamp 1
transform 1 0 34592 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_1174
timestamp 1
transform 1 0 39744 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_1175
timestamp 1
transform 1 0 44896 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_1176
timestamp 1
transform 1 0 50048 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_1177
timestamp 1
transform 1 0 55200 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_1178
timestamp 1
transform 1 0 60352 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_1179
timestamp 1
transform 1 0 65504 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_1180
timestamp 1
transform 1 0 70656 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_1181
timestamp 1
transform 1 0 75808 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_1182
timestamp 1
transform 1 0 80960 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_1183
timestamp 1
transform 1 0 86112 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_1184
timestamp 1
transform 1 0 91264 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_1185
timestamp 1
transform 1 0 96416 0 1 76160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_1186
timestamp 1
transform 1 0 6256 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_1187
timestamp 1
transform 1 0 11408 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_1188
timestamp 1
transform 1 0 16560 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_1189
timestamp 1
transform 1 0 21712 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_1190
timestamp 1
transform 1 0 26864 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_1191
timestamp 1
transform 1 0 32016 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_1192
timestamp 1
transform 1 0 37168 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_1193
timestamp 1
transform 1 0 42320 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_1194
timestamp 1
transform 1 0 47472 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_1195
timestamp 1
transform 1 0 52624 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_1196
timestamp 1
transform 1 0 57776 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_1197
timestamp 1
transform 1 0 62928 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_1198
timestamp 1
transform 1 0 68080 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_1199
timestamp 1
transform 1 0 73232 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_1200
timestamp 1
transform 1 0 78384 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_1201
timestamp 1
transform 1 0 83536 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_1202
timestamp 1
transform 1 0 88688 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_1203
timestamp 1
transform 1 0 93840 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_137_1204
timestamp 1
transform 1 0 98992 0 -1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1205
timestamp 1
transform 1 0 3680 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1206
timestamp 1
transform 1 0 8832 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1207
timestamp 1
transform 1 0 13984 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1208
timestamp 1
transform 1 0 19136 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1209
timestamp 1
transform 1 0 24288 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1210
timestamp 1
transform 1 0 29440 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1211
timestamp 1
transform 1 0 34592 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1212
timestamp 1
transform 1 0 39744 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1213
timestamp 1
transform 1 0 44896 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1214
timestamp 1
transform 1 0 50048 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1215
timestamp 1
transform 1 0 55200 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1216
timestamp 1
transform 1 0 60352 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1217
timestamp 1
transform 1 0 65504 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1218
timestamp 1
transform 1 0 70656 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1219
timestamp 1
transform 1 0 75808 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1220
timestamp 1
transform 1 0 80960 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1221
timestamp 1
transform 1 0 86112 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1222
timestamp 1
transform 1 0 91264 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1223
timestamp 1
transform 1 0 96416 0 1 77248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_139_1224
timestamp 1
transform 1 0 6256 0 -1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_139_1225
timestamp 1
transform 1 0 11408 0 -1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_139_1226
timestamp 1
transform 1 0 16560 0 -1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_139_1227
timestamp 1
transform 1 0 21712 0 -1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_139_1228
timestamp 1
transform 1 0 26864 0 -1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_139_1229
timestamp 1
transform 1 0 32016 0 -1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_139_1230
timestamp 1
transform 1 0 37168 0 -1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_139_1231
timestamp 1
transform 1 0 42320 0 -1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_139_1232
timestamp 1
transform 1 0 47472 0 -1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_139_1233
timestamp 1
transform 1 0 52624 0 -1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_139_1234
timestamp 1
transform 1 0 57776 0 -1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_139_1235
timestamp 1
transform 1 0 62928 0 -1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_139_1236
timestamp 1
transform 1 0 68080 0 -1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_139_1237
timestamp 1
transform 1 0 73232 0 -1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_139_1238
timestamp 1
transform 1 0 78384 0 -1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_139_1239
timestamp 1
transform 1 0 83536 0 -1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_139_1240
timestamp 1
transform 1 0 88688 0 -1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_139_1241
timestamp 1
transform 1 0 93840 0 -1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_139_1242
timestamp 1
transform 1 0 98992 0 -1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_140_1243
timestamp 1
transform 1 0 3680 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_140_1244
timestamp 1
transform 1 0 8832 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_140_1245
timestamp 1
transform 1 0 13984 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_140_1246
timestamp 1
transform 1 0 19136 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_140_1247
timestamp 1
transform 1 0 24288 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_140_1248
timestamp 1
transform 1 0 29440 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_140_1249
timestamp 1
transform 1 0 34592 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_140_1250
timestamp 1
transform 1 0 39744 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_140_1251
timestamp 1
transform 1 0 44896 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_140_1252
timestamp 1
transform 1 0 50048 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_140_1253
timestamp 1
transform 1 0 55200 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_140_1254
timestamp 1
transform 1 0 60352 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_140_1255
timestamp 1
transform 1 0 65504 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_140_1256
timestamp 1
transform 1 0 70656 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_140_1257
timestamp 1
transform 1 0 75808 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_140_1258
timestamp 1
transform 1 0 80960 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_140_1259
timestamp 1
transform 1 0 86112 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_140_1260
timestamp 1
transform 1 0 91264 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_140_1261
timestamp 1
transform 1 0 96416 0 1 78336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_141_1262
timestamp 1
transform 1 0 6256 0 -1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_141_1263
timestamp 1
transform 1 0 11408 0 -1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_141_1264
timestamp 1
transform 1 0 16560 0 -1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_141_1265
timestamp 1
transform 1 0 21712 0 -1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_141_1266
timestamp 1
transform 1 0 26864 0 -1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_141_1267
timestamp 1
transform 1 0 32016 0 -1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_141_1268
timestamp 1
transform 1 0 37168 0 -1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_141_1269
timestamp 1
transform 1 0 42320 0 -1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_141_1270
timestamp 1
transform 1 0 47472 0 -1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_141_1271
timestamp 1
transform 1 0 52624 0 -1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_141_1272
timestamp 1
transform 1 0 57776 0 -1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_141_1273
timestamp 1
transform 1 0 62928 0 -1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_141_1274
timestamp 1
transform 1 0 68080 0 -1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_141_1275
timestamp 1
transform 1 0 73232 0 -1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_141_1276
timestamp 1
transform 1 0 78384 0 -1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_141_1277
timestamp 1
transform 1 0 83536 0 -1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_141_1278
timestamp 1
transform 1 0 88688 0 -1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_141_1279
timestamp 1
transform 1 0 93840 0 -1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_141_1280
timestamp 1
transform 1 0 98992 0 -1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_142_1281
timestamp 1
transform 1 0 3680 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_142_1282
timestamp 1
transform 1 0 8832 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_142_1283
timestamp 1
transform 1 0 13984 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_142_1284
timestamp 1
transform 1 0 19136 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_142_1285
timestamp 1
transform 1 0 24288 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_142_1286
timestamp 1
transform 1 0 29440 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_142_1287
timestamp 1
transform 1 0 34592 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_142_1288
timestamp 1
transform 1 0 39744 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_142_1289
timestamp 1
transform 1 0 44896 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_142_1290
timestamp 1
transform 1 0 50048 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_142_1291
timestamp 1
transform 1 0 55200 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_142_1292
timestamp 1
transform 1 0 60352 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_142_1293
timestamp 1
transform 1 0 65504 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_142_1294
timestamp 1
transform 1 0 70656 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_142_1295
timestamp 1
transform 1 0 75808 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_142_1296
timestamp 1
transform 1 0 80960 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_142_1297
timestamp 1
transform 1 0 86112 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_142_1298
timestamp 1
transform 1 0 91264 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_142_1299
timestamp 1
transform 1 0 96416 0 1 79424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_143_1300
timestamp 1
transform 1 0 6256 0 -1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_143_1301
timestamp 1
transform 1 0 11408 0 -1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_143_1302
timestamp 1
transform 1 0 16560 0 -1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_143_1303
timestamp 1
transform 1 0 21712 0 -1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_143_1304
timestamp 1
transform 1 0 26864 0 -1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_143_1305
timestamp 1
transform 1 0 32016 0 -1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_143_1306
timestamp 1
transform 1 0 37168 0 -1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_143_1307
timestamp 1
transform 1 0 42320 0 -1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_143_1308
timestamp 1
transform 1 0 47472 0 -1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_143_1309
timestamp 1
transform 1 0 52624 0 -1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_143_1310
timestamp 1
transform 1 0 57776 0 -1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_143_1311
timestamp 1
transform 1 0 62928 0 -1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_143_1312
timestamp 1
transform 1 0 68080 0 -1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_143_1313
timestamp 1
transform 1 0 73232 0 -1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_143_1314
timestamp 1
transform 1 0 78384 0 -1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_143_1315
timestamp 1
transform 1 0 83536 0 -1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_143_1316
timestamp 1
transform 1 0 88688 0 -1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_143_1317
timestamp 1
transform 1 0 93840 0 -1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_143_1318
timestamp 1
transform 1 0 98992 0 -1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_144_1319
timestamp 1
transform 1 0 3680 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_144_1320
timestamp 1
transform 1 0 8832 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_144_1321
timestamp 1
transform 1 0 13984 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_144_1322
timestamp 1
transform 1 0 19136 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_144_1323
timestamp 1
transform 1 0 24288 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_144_1324
timestamp 1
transform 1 0 29440 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_144_1325
timestamp 1
transform 1 0 34592 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_144_1326
timestamp 1
transform 1 0 39744 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_144_1327
timestamp 1
transform 1 0 44896 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_144_1328
timestamp 1
transform 1 0 50048 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_144_1329
timestamp 1
transform 1 0 55200 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_144_1330
timestamp 1
transform 1 0 60352 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_144_1331
timestamp 1
transform 1 0 65504 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_144_1332
timestamp 1
transform 1 0 70656 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_144_1333
timestamp 1
transform 1 0 75808 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_144_1334
timestamp 1
transform 1 0 80960 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_144_1335
timestamp 1
transform 1 0 86112 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_144_1336
timestamp 1
transform 1 0 91264 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_144_1337
timestamp 1
transform 1 0 96416 0 1 80512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_145_1338
timestamp 1
transform 1 0 6256 0 -1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_145_1339
timestamp 1
transform 1 0 11408 0 -1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_145_1340
timestamp 1
transform 1 0 16560 0 -1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_145_1341
timestamp 1
transform 1 0 21712 0 -1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_145_1342
timestamp 1
transform 1 0 26864 0 -1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_145_1343
timestamp 1
transform 1 0 32016 0 -1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_145_1344
timestamp 1
transform 1 0 37168 0 -1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_145_1345
timestamp 1
transform 1 0 42320 0 -1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_145_1346
timestamp 1
transform 1 0 47472 0 -1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_145_1347
timestamp 1
transform 1 0 52624 0 -1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_145_1348
timestamp 1
transform 1 0 57776 0 -1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_145_1349
timestamp 1
transform 1 0 62928 0 -1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_145_1350
timestamp 1
transform 1 0 68080 0 -1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_145_1351
timestamp 1
transform 1 0 73232 0 -1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_145_1352
timestamp 1
transform 1 0 78384 0 -1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_145_1353
timestamp 1
transform 1 0 83536 0 -1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_145_1354
timestamp 1
transform 1 0 88688 0 -1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_145_1355
timestamp 1
transform 1 0 93840 0 -1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_145_1356
timestamp 1
transform 1 0 98992 0 -1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_1357
timestamp 1
transform 1 0 3680 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_1358
timestamp 1
transform 1 0 8832 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_1359
timestamp 1
transform 1 0 13984 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_1360
timestamp 1
transform 1 0 19136 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_1361
timestamp 1
transform 1 0 24288 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_1362
timestamp 1
transform 1 0 29440 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_1363
timestamp 1
transform 1 0 34592 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_1364
timestamp 1
transform 1 0 39744 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_1365
timestamp 1
transform 1 0 44896 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_1366
timestamp 1
transform 1 0 50048 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_1367
timestamp 1
transform 1 0 55200 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_1368
timestamp 1
transform 1 0 60352 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_1369
timestamp 1
transform 1 0 65504 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_1370
timestamp 1
transform 1 0 70656 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_1371
timestamp 1
transform 1 0 75808 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_1372
timestamp 1
transform 1 0 80960 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_1373
timestamp 1
transform 1 0 86112 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_1374
timestamp 1
transform 1 0 91264 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_1375
timestamp 1
transform 1 0 96416 0 1 81600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_147_1376
timestamp 1
transform 1 0 6256 0 -1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_147_1377
timestamp 1
transform 1 0 11408 0 -1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_147_1378
timestamp 1
transform 1 0 16560 0 -1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_147_1379
timestamp 1
transform 1 0 21712 0 -1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_147_1380
timestamp 1
transform 1 0 26864 0 -1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_147_1381
timestamp 1
transform 1 0 32016 0 -1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_147_1382
timestamp 1
transform 1 0 37168 0 -1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_147_1383
timestamp 1
transform 1 0 42320 0 -1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_147_1384
timestamp 1
transform 1 0 47472 0 -1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_147_1385
timestamp 1
transform 1 0 52624 0 -1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_147_1386
timestamp 1
transform 1 0 57776 0 -1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_147_1387
timestamp 1
transform 1 0 62928 0 -1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_147_1388
timestamp 1
transform 1 0 68080 0 -1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_147_1389
timestamp 1
transform 1 0 73232 0 -1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_147_1390
timestamp 1
transform 1 0 78384 0 -1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_147_1391
timestamp 1
transform 1 0 83536 0 -1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_147_1392
timestamp 1
transform 1 0 88688 0 -1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_147_1393
timestamp 1
transform 1 0 93840 0 -1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_147_1394
timestamp 1
transform 1 0 98992 0 -1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_1395
timestamp 1
transform 1 0 3680 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_1396
timestamp 1
transform 1 0 8832 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_1397
timestamp 1
transform 1 0 13984 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_1398
timestamp 1
transform 1 0 19136 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_1399
timestamp 1
transform 1 0 24288 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_1400
timestamp 1
transform 1 0 29440 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_1401
timestamp 1
transform 1 0 34592 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_1402
timestamp 1
transform 1 0 39744 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_1403
timestamp 1
transform 1 0 44896 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_1404
timestamp 1
transform 1 0 50048 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_1405
timestamp 1
transform 1 0 55200 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_1406
timestamp 1
transform 1 0 60352 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_1407
timestamp 1
transform 1 0 65504 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_1408
timestamp 1
transform 1 0 70656 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_1409
timestamp 1
transform 1 0 75808 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_1410
timestamp 1
transform 1 0 80960 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_1411
timestamp 1
transform 1 0 86112 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_1412
timestamp 1
transform 1 0 91264 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_1413
timestamp 1
transform 1 0 96416 0 1 82688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_149_1414
timestamp 1
transform 1 0 6256 0 -1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_149_1415
timestamp 1
transform 1 0 11408 0 -1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_149_1416
timestamp 1
transform 1 0 16560 0 -1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_149_1417
timestamp 1
transform 1 0 21712 0 -1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_149_1418
timestamp 1
transform 1 0 26864 0 -1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_149_1419
timestamp 1
transform 1 0 32016 0 -1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_149_1420
timestamp 1
transform 1 0 37168 0 -1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_149_1421
timestamp 1
transform 1 0 42320 0 -1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_149_1422
timestamp 1
transform 1 0 47472 0 -1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_149_1423
timestamp 1
transform 1 0 52624 0 -1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_149_1424
timestamp 1
transform 1 0 57776 0 -1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_149_1425
timestamp 1
transform 1 0 62928 0 -1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_149_1426
timestamp 1
transform 1 0 68080 0 -1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_149_1427
timestamp 1
transform 1 0 73232 0 -1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_149_1428
timestamp 1
transform 1 0 78384 0 -1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_149_1429
timestamp 1
transform 1 0 83536 0 -1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_149_1430
timestamp 1
transform 1 0 88688 0 -1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_149_1431
timestamp 1
transform 1 0 93840 0 -1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_149_1432
timestamp 1
transform 1 0 98992 0 -1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_1433
timestamp 1
transform 1 0 3680 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_1434
timestamp 1
transform 1 0 8832 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_1435
timestamp 1
transform 1 0 13984 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_1436
timestamp 1
transform 1 0 19136 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_1437
timestamp 1
transform 1 0 24288 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_1438
timestamp 1
transform 1 0 29440 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_1439
timestamp 1
transform 1 0 34592 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_1440
timestamp 1
transform 1 0 39744 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_1441
timestamp 1
transform 1 0 44896 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_1442
timestamp 1
transform 1 0 50048 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_1443
timestamp 1
transform 1 0 55200 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_1444
timestamp 1
transform 1 0 60352 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_1445
timestamp 1
transform 1 0 65504 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_1446
timestamp 1
transform 1 0 70656 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_1447
timestamp 1
transform 1 0 75808 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_1448
timestamp 1
transform 1 0 80960 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_1449
timestamp 1
transform 1 0 86112 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_1450
timestamp 1
transform 1 0 91264 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_1451
timestamp 1
transform 1 0 96416 0 1 83776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_1452
timestamp 1
transform 1 0 6256 0 -1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_1453
timestamp 1
transform 1 0 11408 0 -1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_1454
timestamp 1
transform 1 0 16560 0 -1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_1455
timestamp 1
transform 1 0 21712 0 -1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_1456
timestamp 1
transform 1 0 26864 0 -1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_1457
timestamp 1
transform 1 0 32016 0 -1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_1458
timestamp 1
transform 1 0 37168 0 -1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_1459
timestamp 1
transform 1 0 42320 0 -1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_1460
timestamp 1
transform 1 0 47472 0 -1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_1461
timestamp 1
transform 1 0 52624 0 -1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_1462
timestamp 1
transform 1 0 57776 0 -1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_1463
timestamp 1
transform 1 0 62928 0 -1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_1464
timestamp 1
transform 1 0 68080 0 -1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_1465
timestamp 1
transform 1 0 73232 0 -1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_1466
timestamp 1
transform 1 0 78384 0 -1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_1467
timestamp 1
transform 1 0 83536 0 -1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_1468
timestamp 1
transform 1 0 88688 0 -1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_1469
timestamp 1
transform 1 0 93840 0 -1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_1470
timestamp 1
transform 1 0 98992 0 -1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_152_1471
timestamp 1
transform 1 0 3680 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_152_1472
timestamp 1
transform 1 0 8832 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_152_1473
timestamp 1
transform 1 0 13984 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_152_1474
timestamp 1
transform 1 0 19136 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_152_1475
timestamp 1
transform 1 0 24288 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_152_1476
timestamp 1
transform 1 0 29440 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_152_1477
timestamp 1
transform 1 0 34592 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_152_1478
timestamp 1
transform 1 0 39744 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_152_1479
timestamp 1
transform 1 0 44896 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_152_1480
timestamp 1
transform 1 0 50048 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_152_1481
timestamp 1
transform 1 0 55200 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_152_1482
timestamp 1
transform 1 0 60352 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_152_1483
timestamp 1
transform 1 0 65504 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_152_1484
timestamp 1
transform 1 0 70656 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_152_1485
timestamp 1
transform 1 0 75808 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_152_1486
timestamp 1
transform 1 0 80960 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_152_1487
timestamp 1
transform 1 0 86112 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_152_1488
timestamp 1
transform 1 0 91264 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_152_1489
timestamp 1
transform 1 0 96416 0 1 84864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_153_1490
timestamp 1
transform 1 0 6256 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_153_1491
timestamp 1
transform 1 0 11408 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_153_1492
timestamp 1
transform 1 0 16560 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_153_1493
timestamp 1
transform 1 0 21712 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_153_1494
timestamp 1
transform 1 0 26864 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_153_1495
timestamp 1
transform 1 0 32016 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_153_1496
timestamp 1
transform 1 0 37168 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_153_1497
timestamp 1
transform 1 0 42320 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_153_1498
timestamp 1
transform 1 0 47472 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_153_1499
timestamp 1
transform 1 0 52624 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_153_1500
timestamp 1
transform 1 0 57776 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_153_1501
timestamp 1
transform 1 0 62928 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_153_1502
timestamp 1
transform 1 0 68080 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_153_1503
timestamp 1
transform 1 0 73232 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_153_1504
timestamp 1
transform 1 0 78384 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_153_1505
timestamp 1
transform 1 0 83536 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_153_1506
timestamp 1
transform 1 0 88688 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_153_1507
timestamp 1
transform 1 0 93840 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_153_1508
timestamp 1
transform 1 0 98992 0 -1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_1509
timestamp 1
transform 1 0 3680 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_1510
timestamp 1
transform 1 0 8832 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_1511
timestamp 1
transform 1 0 13984 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_1512
timestamp 1
transform 1 0 19136 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_1513
timestamp 1
transform 1 0 24288 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_1514
timestamp 1
transform 1 0 29440 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_1515
timestamp 1
transform 1 0 34592 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_1516
timestamp 1
transform 1 0 39744 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_1517
timestamp 1
transform 1 0 44896 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_1518
timestamp 1
transform 1 0 50048 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_1519
timestamp 1
transform 1 0 55200 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_1520
timestamp 1
transform 1 0 60352 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_1521
timestamp 1
transform 1 0 65504 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_1522
timestamp 1
transform 1 0 70656 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_1523
timestamp 1
transform 1 0 75808 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_1524
timestamp 1
transform 1 0 80960 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_1525
timestamp 1
transform 1 0 86112 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_1526
timestamp 1
transform 1 0 91264 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_1527
timestamp 1
transform 1 0 96416 0 1 85952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_155_1528
timestamp 1
transform 1 0 6256 0 -1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_155_1529
timestamp 1
transform 1 0 11408 0 -1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_155_1530
timestamp 1
transform 1 0 16560 0 -1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_155_1531
timestamp 1
transform 1 0 21712 0 -1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_155_1532
timestamp 1
transform 1 0 26864 0 -1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_155_1533
timestamp 1
transform 1 0 32016 0 -1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_155_1534
timestamp 1
transform 1 0 37168 0 -1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_155_1535
timestamp 1
transform 1 0 42320 0 -1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_155_1536
timestamp 1
transform 1 0 47472 0 -1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_155_1537
timestamp 1
transform 1 0 52624 0 -1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_155_1538
timestamp 1
transform 1 0 57776 0 -1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_155_1539
timestamp 1
transform 1 0 62928 0 -1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_155_1540
timestamp 1
transform 1 0 68080 0 -1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_155_1541
timestamp 1
transform 1 0 73232 0 -1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_155_1542
timestamp 1
transform 1 0 78384 0 -1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_155_1543
timestamp 1
transform 1 0 83536 0 -1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_155_1544
timestamp 1
transform 1 0 88688 0 -1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_155_1545
timestamp 1
transform 1 0 93840 0 -1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_155_1546
timestamp 1
transform 1 0 98992 0 -1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_156_1547
timestamp 1
transform 1 0 3680 0 1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_156_1548
timestamp 1
transform 1 0 8832 0 1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_156_1549
timestamp 1
transform 1 0 13984 0 1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_156_1550
timestamp 1
transform 1 0 19136 0 1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_156_1551
timestamp 1
transform 1 0 24288 0 1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_156_1552
timestamp 1
transform 1 0 29440 0 1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_156_1553
timestamp 1
transform 1 0 34592 0 1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_156_1554
timestamp 1
transform 1 0 39744 0 1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_156_1555
timestamp 1
transform 1 0 44896 0 1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_156_1556
timestamp 1
transform 1 0 50048 0 1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_156_1557
timestamp 1
transform 1 0 55200 0 1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_156_1558
timestamp 1
transform 1 0 60352 0 1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_156_1559
timestamp 1
transform 1 0 65504 0 1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_156_1560
timestamp 1
transform 1 0 70656 0 1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_156_1561
timestamp 1
transform 1 0 75808 0 1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_156_1562
timestamp 1
transform 1 0 80960 0 1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_156_1563
timestamp 1
transform 1 0 86112 0 1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_156_1564
timestamp 1
transform 1 0 91264 0 1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_156_1565
timestamp 1
transform 1 0 96416 0 1 87040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_157_1566
timestamp 1
transform 1 0 6256 0 -1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_157_1567
timestamp 1
transform 1 0 11408 0 -1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_157_1568
timestamp 1
transform 1 0 16560 0 -1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_157_1569
timestamp 1
transform 1 0 21712 0 -1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_157_1570
timestamp 1
transform 1 0 26864 0 -1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_157_1571
timestamp 1
transform 1 0 32016 0 -1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_157_1572
timestamp 1
transform 1 0 37168 0 -1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_157_1573
timestamp 1
transform 1 0 42320 0 -1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_157_1574
timestamp 1
transform 1 0 47472 0 -1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_157_1575
timestamp 1
transform 1 0 52624 0 -1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_157_1576
timestamp 1
transform 1 0 57776 0 -1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_157_1577
timestamp 1
transform 1 0 62928 0 -1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_157_1578
timestamp 1
transform 1 0 68080 0 -1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_157_1579
timestamp 1
transform 1 0 73232 0 -1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_157_1580
timestamp 1
transform 1 0 78384 0 -1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_157_1581
timestamp 1
transform 1 0 83536 0 -1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_157_1582
timestamp 1
transform 1 0 88688 0 -1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_157_1583
timestamp 1
transform 1 0 93840 0 -1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_157_1584
timestamp 1
transform 1 0 98992 0 -1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_158_1585
timestamp 1
transform 1 0 3680 0 1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_158_1586
timestamp 1
transform 1 0 8832 0 1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_158_1587
timestamp 1
transform 1 0 13984 0 1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_158_1588
timestamp 1
transform 1 0 19136 0 1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_158_1589
timestamp 1
transform 1 0 24288 0 1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_158_1590
timestamp 1
transform 1 0 29440 0 1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_158_1591
timestamp 1
transform 1 0 34592 0 1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_158_1592
timestamp 1
transform 1 0 39744 0 1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_158_1593
timestamp 1
transform 1 0 44896 0 1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_158_1594
timestamp 1
transform 1 0 50048 0 1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_158_1595
timestamp 1
transform 1 0 55200 0 1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_158_1596
timestamp 1
transform 1 0 60352 0 1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_158_1597
timestamp 1
transform 1 0 65504 0 1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_158_1598
timestamp 1
transform 1 0 70656 0 1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_158_1599
timestamp 1
transform 1 0 75808 0 1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_158_1600
timestamp 1
transform 1 0 80960 0 1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_158_1601
timestamp 1
transform 1 0 86112 0 1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_158_1602
timestamp 1
transform 1 0 91264 0 1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_158_1603
timestamp 1
transform 1 0 96416 0 1 88128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_159_1604
timestamp 1
transform 1 0 6256 0 -1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_159_1605
timestamp 1
transform 1 0 11408 0 -1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_159_1606
timestamp 1
transform 1 0 16560 0 -1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_159_1607
timestamp 1
transform 1 0 21712 0 -1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_159_1608
timestamp 1
transform 1 0 26864 0 -1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_159_1609
timestamp 1
transform 1 0 32016 0 -1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_159_1610
timestamp 1
transform 1 0 37168 0 -1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_159_1611
timestamp 1
transform 1 0 42320 0 -1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_159_1612
timestamp 1
transform 1 0 47472 0 -1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_159_1613
timestamp 1
transform 1 0 52624 0 -1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_159_1614
timestamp 1
transform 1 0 57776 0 -1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_159_1615
timestamp 1
transform 1 0 62928 0 -1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_159_1616
timestamp 1
transform 1 0 68080 0 -1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_159_1617
timestamp 1
transform 1 0 73232 0 -1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_159_1618
timestamp 1
transform 1 0 78384 0 -1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_159_1619
timestamp 1
transform 1 0 83536 0 -1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_159_1620
timestamp 1
transform 1 0 88688 0 -1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_159_1621
timestamp 1
transform 1 0 93840 0 -1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_159_1622
timestamp 1
transform 1 0 98992 0 -1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_160_1623
timestamp 1
transform 1 0 3680 0 1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_160_1624
timestamp 1
transform 1 0 8832 0 1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_160_1625
timestamp 1
transform 1 0 13984 0 1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_160_1626
timestamp 1
transform 1 0 19136 0 1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_160_1627
timestamp 1
transform 1 0 24288 0 1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_160_1628
timestamp 1
transform 1 0 29440 0 1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_160_1629
timestamp 1
transform 1 0 34592 0 1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_160_1630
timestamp 1
transform 1 0 39744 0 1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_160_1631
timestamp 1
transform 1 0 44896 0 1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_160_1632
timestamp 1
transform 1 0 50048 0 1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_160_1633
timestamp 1
transform 1 0 55200 0 1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_160_1634
timestamp 1
transform 1 0 60352 0 1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_160_1635
timestamp 1
transform 1 0 65504 0 1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_160_1636
timestamp 1
transform 1 0 70656 0 1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_160_1637
timestamp 1
transform 1 0 75808 0 1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_160_1638
timestamp 1
transform 1 0 80960 0 1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_160_1639
timestamp 1
transform 1 0 86112 0 1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_160_1640
timestamp 1
transform 1 0 91264 0 1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_160_1641
timestamp 1
transform 1 0 96416 0 1 89216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_161_1642
timestamp 1
transform 1 0 6256 0 -1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_161_1643
timestamp 1
transform 1 0 11408 0 -1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_161_1644
timestamp 1
transform 1 0 16560 0 -1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_161_1645
timestamp 1
transform 1 0 21712 0 -1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_161_1646
timestamp 1
transform 1 0 26864 0 -1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_161_1647
timestamp 1
transform 1 0 32016 0 -1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_161_1648
timestamp 1
transform 1 0 37168 0 -1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_161_1649
timestamp 1
transform 1 0 42320 0 -1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_161_1650
timestamp 1
transform 1 0 47472 0 -1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_161_1651
timestamp 1
transform 1 0 52624 0 -1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_161_1652
timestamp 1
transform 1 0 57776 0 -1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_161_1653
timestamp 1
transform 1 0 62928 0 -1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_161_1654
timestamp 1
transform 1 0 68080 0 -1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_161_1655
timestamp 1
transform 1 0 73232 0 -1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_161_1656
timestamp 1
transform 1 0 78384 0 -1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_161_1657
timestamp 1
transform 1 0 83536 0 -1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_161_1658
timestamp 1
transform 1 0 88688 0 -1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_161_1659
timestamp 1
transform 1 0 93840 0 -1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_161_1660
timestamp 1
transform 1 0 98992 0 -1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_162_1661
timestamp 1
transform 1 0 3680 0 1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_162_1662
timestamp 1
transform 1 0 8832 0 1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_162_1663
timestamp 1
transform 1 0 13984 0 1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_162_1664
timestamp 1
transform 1 0 19136 0 1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_162_1665
timestamp 1
transform 1 0 24288 0 1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_162_1666
timestamp 1
transform 1 0 29440 0 1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_162_1667
timestamp 1
transform 1 0 34592 0 1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_162_1668
timestamp 1
transform 1 0 39744 0 1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_162_1669
timestamp 1
transform 1 0 44896 0 1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_162_1670
timestamp 1
transform 1 0 50048 0 1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_162_1671
timestamp 1
transform 1 0 55200 0 1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_162_1672
timestamp 1
transform 1 0 60352 0 1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_162_1673
timestamp 1
transform 1 0 65504 0 1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_162_1674
timestamp 1
transform 1 0 70656 0 1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_162_1675
timestamp 1
transform 1 0 75808 0 1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_162_1676
timestamp 1
transform 1 0 80960 0 1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_162_1677
timestamp 1
transform 1 0 86112 0 1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_162_1678
timestamp 1
transform 1 0 91264 0 1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_162_1679
timestamp 1
transform 1 0 96416 0 1 90304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_163_1680
timestamp 1
transform 1 0 6256 0 -1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_163_1681
timestamp 1
transform 1 0 11408 0 -1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_163_1682
timestamp 1
transform 1 0 16560 0 -1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_163_1683
timestamp 1
transform 1 0 21712 0 -1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_163_1684
timestamp 1
transform 1 0 26864 0 -1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_163_1685
timestamp 1
transform 1 0 32016 0 -1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_163_1686
timestamp 1
transform 1 0 37168 0 -1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_163_1687
timestamp 1
transform 1 0 42320 0 -1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_163_1688
timestamp 1
transform 1 0 47472 0 -1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_163_1689
timestamp 1
transform 1 0 52624 0 -1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_163_1690
timestamp 1
transform 1 0 57776 0 -1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_163_1691
timestamp 1
transform 1 0 62928 0 -1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_163_1692
timestamp 1
transform 1 0 68080 0 -1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_163_1693
timestamp 1
transform 1 0 73232 0 -1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_163_1694
timestamp 1
transform 1 0 78384 0 -1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_163_1695
timestamp 1
transform 1 0 83536 0 -1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_163_1696
timestamp 1
transform 1 0 88688 0 -1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_163_1697
timestamp 1
transform 1 0 93840 0 -1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_163_1698
timestamp 1
transform 1 0 98992 0 -1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_164_1699
timestamp 1
transform 1 0 3680 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_164_1700
timestamp 1
transform 1 0 8832 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_164_1701
timestamp 1
transform 1 0 13984 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_164_1702
timestamp 1
transform 1 0 19136 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_164_1703
timestamp 1
transform 1 0 24288 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_164_1704
timestamp 1
transform 1 0 29440 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_164_1705
timestamp 1
transform 1 0 34592 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_164_1706
timestamp 1
transform 1 0 39744 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_164_1707
timestamp 1
transform 1 0 44896 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_164_1708
timestamp 1
transform 1 0 50048 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_164_1709
timestamp 1
transform 1 0 55200 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_164_1710
timestamp 1
transform 1 0 60352 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_164_1711
timestamp 1
transform 1 0 65504 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_164_1712
timestamp 1
transform 1 0 70656 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_164_1713
timestamp 1
transform 1 0 75808 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_164_1714
timestamp 1
transform 1 0 80960 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_164_1715
timestamp 1
transform 1 0 86112 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_164_1716
timestamp 1
transform 1 0 91264 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_164_1717
timestamp 1
transform 1 0 96416 0 1 91392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_1718
timestamp 1
transform 1 0 6256 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_1719
timestamp 1
transform 1 0 11408 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_1720
timestamp 1
transform 1 0 16560 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_1721
timestamp 1
transform 1 0 21712 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_1722
timestamp 1
transform 1 0 26864 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_1723
timestamp 1
transform 1 0 32016 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_1724
timestamp 1
transform 1 0 37168 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_1725
timestamp 1
transform 1 0 42320 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_1726
timestamp 1
transform 1 0 47472 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_1727
timestamp 1
transform 1 0 52624 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_1728
timestamp 1
transform 1 0 57776 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_1729
timestamp 1
transform 1 0 62928 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_1730
timestamp 1
transform 1 0 68080 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_1731
timestamp 1
transform 1 0 73232 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_1732
timestamp 1
transform 1 0 78384 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_1733
timestamp 1
transform 1 0 83536 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_1734
timestamp 1
transform 1 0 88688 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_1735
timestamp 1
transform 1 0 93840 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_165_1736
timestamp 1
transform 1 0 98992 0 -1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_166_1737
timestamp 1
transform 1 0 3680 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_166_1738
timestamp 1
transform 1 0 8832 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_166_1739
timestamp 1
transform 1 0 13984 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_166_1740
timestamp 1
transform 1 0 19136 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_166_1741
timestamp 1
transform 1 0 24288 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_166_1742
timestamp 1
transform 1 0 29440 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_166_1743
timestamp 1
transform 1 0 34592 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_166_1744
timestamp 1
transform 1 0 39744 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_166_1745
timestamp 1
transform 1 0 44896 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_166_1746
timestamp 1
transform 1 0 50048 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_166_1747
timestamp 1
transform 1 0 55200 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_166_1748
timestamp 1
transform 1 0 60352 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_166_1749
timestamp 1
transform 1 0 65504 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_166_1750
timestamp 1
transform 1 0 70656 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_166_1751
timestamp 1
transform 1 0 75808 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_166_1752
timestamp 1
transform 1 0 80960 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_166_1753
timestamp 1
transform 1 0 86112 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_166_1754
timestamp 1
transform 1 0 91264 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_166_1755
timestamp 1
transform 1 0 96416 0 1 92480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_1756
timestamp 1
transform 1 0 6256 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_1757
timestamp 1
transform 1 0 11408 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_1758
timestamp 1
transform 1 0 16560 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_1759
timestamp 1
transform 1 0 21712 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_1760
timestamp 1
transform 1 0 26864 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_1761
timestamp 1
transform 1 0 32016 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_1762
timestamp 1
transform 1 0 37168 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_1763
timestamp 1
transform 1 0 42320 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_1764
timestamp 1
transform 1 0 47472 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_1765
timestamp 1
transform 1 0 52624 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_1766
timestamp 1
transform 1 0 57776 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_1767
timestamp 1
transform 1 0 62928 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_1768
timestamp 1
transform 1 0 68080 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_1769
timestamp 1
transform 1 0 73232 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_1770
timestamp 1
transform 1 0 78384 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_1771
timestamp 1
transform 1 0 83536 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_1772
timestamp 1
transform 1 0 88688 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_1773
timestamp 1
transform 1 0 93840 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_167_1774
timestamp 1
transform 1 0 98992 0 -1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_1775
timestamp 1
transform 1 0 3680 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_1776
timestamp 1
transform 1 0 8832 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_1777
timestamp 1
transform 1 0 13984 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_1778
timestamp 1
transform 1 0 19136 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_1779
timestamp 1
transform 1 0 24288 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_1780
timestamp 1
transform 1 0 29440 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_1781
timestamp 1
transform 1 0 34592 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_1782
timestamp 1
transform 1 0 39744 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_1783
timestamp 1
transform 1 0 44896 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_1784
timestamp 1
transform 1 0 50048 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_1785
timestamp 1
transform 1 0 55200 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_1786
timestamp 1
transform 1 0 60352 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_1787
timestamp 1
transform 1 0 65504 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_1788
timestamp 1
transform 1 0 70656 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_1789
timestamp 1
transform 1 0 75808 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_1790
timestamp 1
transform 1 0 80960 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_1791
timestamp 1
transform 1 0 86112 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_1792
timestamp 1
transform 1 0 91264 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_168_1793
timestamp 1
transform 1 0 96416 0 1 93568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_1794
timestamp 1
transform 1 0 6256 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_1795
timestamp 1
transform 1 0 11408 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_1796
timestamp 1
transform 1 0 16560 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_1797
timestamp 1
transform 1 0 21712 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_1798
timestamp 1
transform 1 0 26864 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_1799
timestamp 1
transform 1 0 32016 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_1800
timestamp 1
transform 1 0 37168 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_1801
timestamp 1
transform 1 0 42320 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_1802
timestamp 1
transform 1 0 47472 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_1803
timestamp 1
transform 1 0 52624 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_1804
timestamp 1
transform 1 0 57776 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_1805
timestamp 1
transform 1 0 62928 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_1806
timestamp 1
transform 1 0 68080 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_1807
timestamp 1
transform 1 0 73232 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_1808
timestamp 1
transform 1 0 78384 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_1809
timestamp 1
transform 1 0 83536 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_1810
timestamp 1
transform 1 0 88688 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_1811
timestamp 1
transform 1 0 93840 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_169_1812
timestamp 1
transform 1 0 98992 0 -1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_1813
timestamp 1
transform 1 0 3680 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_1814
timestamp 1
transform 1 0 8832 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_1815
timestamp 1
transform 1 0 13984 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_1816
timestamp 1
transform 1 0 19136 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_1817
timestamp 1
transform 1 0 24288 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_1818
timestamp 1
transform 1 0 29440 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_1819
timestamp 1
transform 1 0 34592 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_1820
timestamp 1
transform 1 0 39744 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_1821
timestamp 1
transform 1 0 44896 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_1822
timestamp 1
transform 1 0 50048 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_1823
timestamp 1
transform 1 0 55200 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_1824
timestamp 1
transform 1 0 60352 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_1825
timestamp 1
transform 1 0 65504 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_1826
timestamp 1
transform 1 0 70656 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_1827
timestamp 1
transform 1 0 75808 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_1828
timestamp 1
transform 1 0 80960 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_1829
timestamp 1
transform 1 0 86112 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_1830
timestamp 1
transform 1 0 91264 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_170_1831
timestamp 1
transform 1 0 96416 0 1 94656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1832
timestamp 1
transform 1 0 6256 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1833
timestamp 1
transform 1 0 11408 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1834
timestamp 1
transform 1 0 16560 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1835
timestamp 1
transform 1 0 21712 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1836
timestamp 1
transform 1 0 26864 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1837
timestamp 1
transform 1 0 32016 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1838
timestamp 1
transform 1 0 37168 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1839
timestamp 1
transform 1 0 42320 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1840
timestamp 1
transform 1 0 47472 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1841
timestamp 1
transform 1 0 52624 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1842
timestamp 1
transform 1 0 57776 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1843
timestamp 1
transform 1 0 62928 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1844
timestamp 1
transform 1 0 68080 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1845
timestamp 1
transform 1 0 73232 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1846
timestamp 1
transform 1 0 78384 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1847
timestamp 1
transform 1 0 83536 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1848
timestamp 1
transform 1 0 88688 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1849
timestamp 1
transform 1 0 93840 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_171_1850
timestamp 1
transform 1 0 98992 0 -1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_172_1851
timestamp 1
transform 1 0 3680 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_172_1852
timestamp 1
transform 1 0 8832 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_172_1853
timestamp 1
transform 1 0 13984 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_172_1854
timestamp 1
transform 1 0 19136 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_172_1855
timestamp 1
transform 1 0 24288 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_172_1856
timestamp 1
transform 1 0 29440 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_172_1857
timestamp 1
transform 1 0 34592 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_172_1858
timestamp 1
transform 1 0 39744 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_172_1859
timestamp 1
transform 1 0 44896 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_172_1860
timestamp 1
transform 1 0 50048 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_172_1861
timestamp 1
transform 1 0 55200 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_172_1862
timestamp 1
transform 1 0 60352 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_172_1863
timestamp 1
transform 1 0 65504 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_172_1864
timestamp 1
transform 1 0 70656 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_172_1865
timestamp 1
transform 1 0 75808 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_172_1866
timestamp 1
transform 1 0 80960 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_172_1867
timestamp 1
transform 1 0 86112 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_172_1868
timestamp 1
transform 1 0 91264 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_172_1869
timestamp 1
transform 1 0 96416 0 1 95744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_173_1870
timestamp 1
transform 1 0 6256 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_173_1871
timestamp 1
transform 1 0 11408 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_173_1872
timestamp 1
transform 1 0 16560 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_173_1873
timestamp 1
transform 1 0 21712 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_173_1874
timestamp 1
transform 1 0 26864 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_173_1875
timestamp 1
transform 1 0 32016 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_173_1876
timestamp 1
transform 1 0 37168 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_173_1877
timestamp 1
transform 1 0 42320 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_173_1878
timestamp 1
transform 1 0 47472 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_173_1879
timestamp 1
transform 1 0 52624 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_173_1880
timestamp 1
transform 1 0 57776 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_173_1881
timestamp 1
transform 1 0 62928 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_173_1882
timestamp 1
transform 1 0 68080 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_173_1883
timestamp 1
transform 1 0 73232 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_173_1884
timestamp 1
transform 1 0 78384 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_173_1885
timestamp 1
transform 1 0 83536 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_173_1886
timestamp 1
transform 1 0 88688 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_173_1887
timestamp 1
transform 1 0 93840 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_173_1888
timestamp 1
transform 1 0 98992 0 -1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_1889
timestamp 1
transform 1 0 3680 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_1890
timestamp 1
transform 1 0 8832 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_1891
timestamp 1
transform 1 0 13984 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_1892
timestamp 1
transform 1 0 19136 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_1893
timestamp 1
transform 1 0 24288 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_1894
timestamp 1
transform 1 0 29440 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_1895
timestamp 1
transform 1 0 34592 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_1896
timestamp 1
transform 1 0 39744 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_1897
timestamp 1
transform 1 0 44896 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_1898
timestamp 1
transform 1 0 50048 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_1899
timestamp 1
transform 1 0 55200 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_1900
timestamp 1
transform 1 0 60352 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_1901
timestamp 1
transform 1 0 65504 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_1902
timestamp 1
transform 1 0 70656 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_1903
timestamp 1
transform 1 0 75808 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_1904
timestamp 1
transform 1 0 80960 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_1905
timestamp 1
transform 1 0 86112 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_1906
timestamp 1
transform 1 0 91264 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_174_1907
timestamp 1
transform 1 0 96416 0 1 96832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_175_1908
timestamp 1
transform 1 0 6256 0 -1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_175_1909
timestamp 1
transform 1 0 11408 0 -1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_175_1910
timestamp 1
transform 1 0 16560 0 -1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_175_1911
timestamp 1
transform 1 0 21712 0 -1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_175_1912
timestamp 1
transform 1 0 26864 0 -1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_175_1913
timestamp 1
transform 1 0 32016 0 -1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_175_1914
timestamp 1
transform 1 0 37168 0 -1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_175_1915
timestamp 1
transform 1 0 42320 0 -1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_175_1916
timestamp 1
transform 1 0 47472 0 -1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_175_1917
timestamp 1
transform 1 0 52624 0 -1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_175_1918
timestamp 1
transform 1 0 57776 0 -1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_175_1919
timestamp 1
transform 1 0 62928 0 -1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_175_1920
timestamp 1
transform 1 0 68080 0 -1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_175_1921
timestamp 1
transform 1 0 73232 0 -1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_175_1922
timestamp 1
transform 1 0 78384 0 -1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_175_1923
timestamp 1
transform 1 0 83536 0 -1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_175_1924
timestamp 1
transform 1 0 88688 0 -1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_175_1925
timestamp 1
transform 1 0 93840 0 -1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_175_1926
timestamp 1
transform 1 0 98992 0 -1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_176_1927
timestamp 1
transform 1 0 3680 0 1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_176_1928
timestamp 1
transform 1 0 8832 0 1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_176_1929
timestamp 1
transform 1 0 13984 0 1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_176_1930
timestamp 1
transform 1 0 19136 0 1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_176_1931
timestamp 1
transform 1 0 24288 0 1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_176_1932
timestamp 1
transform 1 0 29440 0 1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_176_1933
timestamp 1
transform 1 0 34592 0 1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_176_1934
timestamp 1
transform 1 0 39744 0 1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_176_1935
timestamp 1
transform 1 0 44896 0 1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_176_1936
timestamp 1
transform 1 0 50048 0 1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_176_1937
timestamp 1
transform 1 0 55200 0 1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_176_1938
timestamp 1
transform 1 0 60352 0 1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_176_1939
timestamp 1
transform 1 0 65504 0 1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_176_1940
timestamp 1
transform 1 0 70656 0 1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_176_1941
timestamp 1
transform 1 0 75808 0 1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_176_1942
timestamp 1
transform 1 0 80960 0 1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_176_1943
timestamp 1
transform 1 0 86112 0 1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_176_1944
timestamp 1
transform 1 0 91264 0 1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_176_1945
timestamp 1
transform 1 0 96416 0 1 97920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_177_1946
timestamp 1
transform 1 0 6256 0 -1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_177_1947
timestamp 1
transform 1 0 11408 0 -1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_177_1948
timestamp 1
transform 1 0 16560 0 -1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_177_1949
timestamp 1
transform 1 0 21712 0 -1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_177_1950
timestamp 1
transform 1 0 26864 0 -1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_177_1951
timestamp 1
transform 1 0 32016 0 -1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_177_1952
timestamp 1
transform 1 0 37168 0 -1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_177_1953
timestamp 1
transform 1 0 42320 0 -1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_177_1954
timestamp 1
transform 1 0 47472 0 -1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_177_1955
timestamp 1
transform 1 0 52624 0 -1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_177_1956
timestamp 1
transform 1 0 57776 0 -1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_177_1957
timestamp 1
transform 1 0 62928 0 -1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_177_1958
timestamp 1
transform 1 0 68080 0 -1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_177_1959
timestamp 1
transform 1 0 73232 0 -1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_177_1960
timestamp 1
transform 1 0 78384 0 -1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_177_1961
timestamp 1
transform 1 0 83536 0 -1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_177_1962
timestamp 1
transform 1 0 88688 0 -1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_177_1963
timestamp 1
transform 1 0 93840 0 -1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_177_1964
timestamp 1
transform 1 0 98992 0 -1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_178_1965
timestamp 1
transform 1 0 3680 0 1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_178_1966
timestamp 1
transform 1 0 8832 0 1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_178_1967
timestamp 1
transform 1 0 13984 0 1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_178_1968
timestamp 1
transform 1 0 19136 0 1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_178_1969
timestamp 1
transform 1 0 24288 0 1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_178_1970
timestamp 1
transform 1 0 29440 0 1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_178_1971
timestamp 1
transform 1 0 34592 0 1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_178_1972
timestamp 1
transform 1 0 39744 0 1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_178_1973
timestamp 1
transform 1 0 44896 0 1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_178_1974
timestamp 1
transform 1 0 50048 0 1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_178_1975
timestamp 1
transform 1 0 55200 0 1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_178_1976
timestamp 1
transform 1 0 60352 0 1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_178_1977
timestamp 1
transform 1 0 65504 0 1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_178_1978
timestamp 1
transform 1 0 70656 0 1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_178_1979
timestamp 1
transform 1 0 75808 0 1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_178_1980
timestamp 1
transform 1 0 80960 0 1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_178_1981
timestamp 1
transform 1 0 86112 0 1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_178_1982
timestamp 1
transform 1 0 91264 0 1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_178_1983
timestamp 1
transform 1 0 96416 0 1 99008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_179_1984
timestamp 1
transform 1 0 6256 0 -1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_179_1985
timestamp 1
transform 1 0 11408 0 -1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_179_1986
timestamp 1
transform 1 0 16560 0 -1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_179_1987
timestamp 1
transform 1 0 21712 0 -1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_179_1988
timestamp 1
transform 1 0 26864 0 -1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_179_1989
timestamp 1
transform 1 0 32016 0 -1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_179_1990
timestamp 1
transform 1 0 37168 0 -1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_179_1991
timestamp 1
transform 1 0 42320 0 -1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_179_1992
timestamp 1
transform 1 0 47472 0 -1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_179_1993
timestamp 1
transform 1 0 52624 0 -1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_179_1994
timestamp 1
transform 1 0 57776 0 -1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_179_1995
timestamp 1
transform 1 0 62928 0 -1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_179_1996
timestamp 1
transform 1 0 68080 0 -1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_179_1997
timestamp 1
transform 1 0 73232 0 -1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_179_1998
timestamp 1
transform 1 0 78384 0 -1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_179_1999
timestamp 1
transform 1 0 83536 0 -1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_179_2000
timestamp 1
transform 1 0 88688 0 -1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_179_2001
timestamp 1
transform 1 0 93840 0 -1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_179_2002
timestamp 1
transform 1 0 98992 0 -1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_180_2003
timestamp 1
transform 1 0 3680 0 1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_180_2004
timestamp 1
transform 1 0 8832 0 1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_180_2005
timestamp 1
transform 1 0 13984 0 1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_180_2006
timestamp 1
transform 1 0 19136 0 1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_180_2007
timestamp 1
transform 1 0 24288 0 1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_180_2008
timestamp 1
transform 1 0 29440 0 1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_180_2009
timestamp 1
transform 1 0 34592 0 1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_180_2010
timestamp 1
transform 1 0 39744 0 1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_180_2011
timestamp 1
transform 1 0 44896 0 1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_180_2012
timestamp 1
transform 1 0 50048 0 1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_180_2013
timestamp 1
transform 1 0 55200 0 1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_180_2014
timestamp 1
transform 1 0 60352 0 1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_180_2015
timestamp 1
transform 1 0 65504 0 1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_180_2016
timestamp 1
transform 1 0 70656 0 1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_180_2017
timestamp 1
transform 1 0 75808 0 1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_180_2018
timestamp 1
transform 1 0 80960 0 1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_180_2019
timestamp 1
transform 1 0 86112 0 1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_180_2020
timestamp 1
transform 1 0 91264 0 1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_180_2021
timestamp 1
transform 1 0 96416 0 1 100096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_181_2022
timestamp 1
transform 1 0 6256 0 -1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_181_2023
timestamp 1
transform 1 0 11408 0 -1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_181_2024
timestamp 1
transform 1 0 16560 0 -1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_181_2025
timestamp 1
transform 1 0 21712 0 -1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_181_2026
timestamp 1
transform 1 0 26864 0 -1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_181_2027
timestamp 1
transform 1 0 32016 0 -1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_181_2028
timestamp 1
transform 1 0 37168 0 -1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_181_2029
timestamp 1
transform 1 0 42320 0 -1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_181_2030
timestamp 1
transform 1 0 47472 0 -1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_181_2031
timestamp 1
transform 1 0 52624 0 -1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_181_2032
timestamp 1
transform 1 0 57776 0 -1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_181_2033
timestamp 1
transform 1 0 62928 0 -1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_181_2034
timestamp 1
transform 1 0 68080 0 -1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_181_2035
timestamp 1
transform 1 0 73232 0 -1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_181_2036
timestamp 1
transform 1 0 78384 0 -1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_181_2037
timestamp 1
transform 1 0 83536 0 -1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_181_2038
timestamp 1
transform 1 0 88688 0 -1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_181_2039
timestamp 1
transform 1 0 93840 0 -1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_181_2040
timestamp 1
transform 1 0 98992 0 -1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_182_2041
timestamp 1
transform 1 0 3680 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_182_2042
timestamp 1
transform 1 0 6256 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_182_2043
timestamp 1
transform 1 0 8832 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_182_2044
timestamp 1
transform 1 0 11408 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_182_2045
timestamp 1
transform 1 0 13984 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_182_2046
timestamp 1
transform 1 0 16560 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_182_2047
timestamp 1
transform 1 0 19136 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_182_2048
timestamp 1
transform 1 0 21712 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_182_2049
timestamp 1
transform 1 0 24288 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_182_2050
timestamp 1
transform 1 0 26864 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_182_2051
timestamp 1
transform 1 0 29440 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_182_2052
timestamp 1
transform 1 0 32016 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_182_2053
timestamp 1
transform 1 0 34592 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_182_2054
timestamp 1
transform 1 0 37168 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_182_2055
timestamp 1
transform 1 0 39744 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_182_2056
timestamp 1
transform 1 0 42320 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_182_2057
timestamp 1
transform 1 0 44896 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_182_2058
timestamp 1
transform 1 0 47472 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_182_2059
timestamp 1
transform 1 0 50048 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_182_2060
timestamp 1
transform 1 0 52624 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_182_2061
timestamp 1
transform 1 0 55200 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_182_2062
timestamp 1
transform 1 0 57776 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_182_2063
timestamp 1
transform 1 0 60352 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_182_2064
timestamp 1
transform 1 0 62928 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_182_2065
timestamp 1
transform 1 0 65504 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_182_2066
timestamp 1
transform 1 0 68080 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_182_2067
timestamp 1
transform 1 0 70656 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_182_2068
timestamp 1
transform 1 0 73232 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_182_2069
timestamp 1
transform 1 0 75808 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_182_2070
timestamp 1
transform 1 0 78384 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_182_2071
timestamp 1
transform 1 0 80960 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_182_2072
timestamp 1
transform 1 0 83536 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_182_2073
timestamp 1
transform 1 0 86112 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_182_2074
timestamp 1
transform 1 0 88688 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_182_2075
timestamp 1
transform 1 0 91264 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_182_2076
timestamp 1
transform 1 0 93840 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_182_2077
timestamp 1
transform 1 0 96416 0 1 101184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_182_2078
timestamp 1
transform 1 0 98992 0 1 101184
box -38 -48 130 592
<< labels >>
flabel metal2 s 17406 0 17462 800 0 FreeSans 224 90 0 0 addr0[0]
port 0 nsew signal input
flabel metal2 s 18694 0 18750 800 0 FreeSans 224 90 0 0 addr0[1]
port 1 nsew signal input
flabel metal3 s 0 27888 800 28008 0 FreeSans 480 0 0 0 addr0[2]
port 2 nsew signal input
flabel metal3 s 0 29248 800 29368 0 FreeSans 480 0 0 0 addr0[3]
port 3 nsew signal input
flabel metal3 s 0 30608 800 30728 0 FreeSans 480 0 0 0 addr0[4]
port 4 nsew signal input
flabel metal3 s 0 32648 800 32768 0 FreeSans 480 0 0 0 addr0[5]
port 5 nsew signal input
flabel metal3 s 0 33328 800 33448 0 FreeSans 480 0 0 0 addr0[6]
port 6 nsew signal input
flabel metal3 s 0 35368 800 35488 0 FreeSans 480 0 0 0 addr0[7]
port 7 nsew signal input
flabel metal3 s 101162 4088 101962 4208 0 FreeSans 480 0 0 0 clk
port 8 nsew signal input
flabel metal3 s 0 9528 800 9648 0 FreeSans 480 0 0 0 csb0
port 9 nsew signal input
flabel metal2 s 19982 0 20038 800 0 FreeSans 224 90 0 0 din0[0]
port 10 nsew signal input
flabel metal2 s 31574 0 31630 800 0 FreeSans 224 90 0 0 din0[10]
port 11 nsew signal input
flabel metal2 s 32862 0 32918 800 0 FreeSans 224 90 0 0 din0[11]
port 12 nsew signal input
flabel metal2 s 33506 0 33562 800 0 FreeSans 224 90 0 0 din0[12]
port 13 nsew signal input
flabel metal2 s 34794 0 34850 800 0 FreeSans 224 90 0 0 din0[13]
port 14 nsew signal input
flabel metal2 s 36082 0 36138 800 0 FreeSans 224 90 0 0 din0[14]
port 15 nsew signal input
flabel metal2 s 37370 0 37426 800 0 FreeSans 224 90 0 0 din0[15]
port 16 nsew signal input
flabel metal2 s 20626 0 20682 800 0 FreeSans 224 90 0 0 din0[1]
port 17 nsew signal input
flabel metal2 s 21914 0 21970 800 0 FreeSans 224 90 0 0 din0[2]
port 18 nsew signal input
flabel metal2 s 23202 0 23258 800 0 FreeSans 224 90 0 0 din0[3]
port 19 nsew signal input
flabel metal2 s 24490 0 24546 800 0 FreeSans 224 90 0 0 din0[4]
port 20 nsew signal input
flabel metal2 s 25778 0 25834 800 0 FreeSans 224 90 0 0 din0[5]
port 21 nsew signal input
flabel metal2 s 27066 0 27122 800 0 FreeSans 224 90 0 0 din0[6]
port 22 nsew signal input
flabel metal2 s 27710 0 27766 800 0 FreeSans 224 90 0 0 din0[7]
port 23 nsew signal input
flabel metal2 s 28998 0 29054 800 0 FreeSans 224 90 0 0 din0[8]
port 24 nsew signal input
flabel metal2 s 30286 0 30342 800 0 FreeSans 224 90 0 0 din0[9]
port 25 nsew signal input
flabel metal3 s 101162 25848 101962 25968 0 FreeSans 480 0 0 0 rst
port 26 nsew signal input
flabel metal3 s 0 61208 800 61328 0 FreeSans 480 0 0 0 sine_out[0]
port 27 nsew signal output
flabel metal2 s 58622 103306 58678 104106 0 FreeSans 224 90 0 0 sine_out[10]
port 28 nsew signal output
flabel metal3 s 101162 62568 101962 62688 0 FreeSans 480 0 0 0 sine_out[11]
port 29 nsew signal output
flabel metal3 s 101162 61888 101962 62008 0 FreeSans 480 0 0 0 sine_out[12]
port 30 nsew signal output
flabel metal3 s 101162 59848 101962 59968 0 FreeSans 480 0 0 0 sine_out[13]
port 31 nsew signal output
flabel metal3 s 101162 61208 101962 61328 0 FreeSans 480 0 0 0 sine_out[14]
port 32 nsew signal output
flabel metal3 s 101162 60528 101962 60648 0 FreeSans 480 0 0 0 sine_out[15]
port 33 nsew signal output
flabel metal3 s 0 61888 800 62008 0 FreeSans 480 0 0 0 sine_out[1]
port 34 nsew signal output
flabel metal2 s 43166 103306 43222 104106 0 FreeSans 224 90 0 0 sine_out[2]
port 35 nsew signal output
flabel metal2 s 45098 103306 45154 104106 0 FreeSans 224 90 0 0 sine_out[3]
port 36 nsew signal output
flabel metal2 s 47674 103306 47730 104106 0 FreeSans 224 90 0 0 sine_out[4]
port 37 nsew signal output
flabel metal2 s 49606 103306 49662 104106 0 FreeSans 224 90 0 0 sine_out[5]
port 38 nsew signal output
flabel metal2 s 50894 103306 50950 104106 0 FreeSans 224 90 0 0 sine_out[6]
port 39 nsew signal output
flabel metal2 s 52826 103306 52882 104106 0 FreeSans 224 90 0 0 sine_out[7]
port 40 nsew signal output
flabel metal2 s 55402 103306 55458 104106 0 FreeSans 224 90 0 0 sine_out[8]
port 41 nsew signal output
flabel metal2 s 57334 103306 57390 104106 0 FreeSans 224 90 0 0 sine_out[9]
port 42 nsew signal output
flabel metal4 s 4208 59834 4528 101776 0 FreeSans 1920 90 0 0 vccd1
port 43 nsew power bidirectional
flabel metal4 s 34928 59834 35248 101776 0 FreeSans 1920 90 0 0 vccd1
port 43 nsew power bidirectional
flabel metal4 s 65648 59650 65968 101776 0 FreeSans 1920 90 0 0 vccd1
port 43 nsew power bidirectional
flabel metal4 s 96368 59650 96688 101776 0 FreeSans 1920 90 0 0 vccd1
port 43 nsew power bidirectional
flabel metal5 s 1056 5346 100880 5666 0 FreeSans 2560 0 0 0 vccd1
port 43 nsew power bidirectional
flabel metal5 s 1056 35982 100880 36302 0 FreeSans 2560 0 0 0 vccd1
port 43 nsew power bidirectional
flabel metal5 s 1056 66618 100880 66938 0 FreeSans 2560 0 0 0 vccd1
port 43 nsew power bidirectional
flabel metal5 s 1056 97254 100880 97574 0 FreeSans 2560 0 0 0 vccd1
port 43 nsew power bidirectional
flabel metal4 s 1300 2128 1460 60432 0 FreeSans 960 90 0 0 vccd1
port 43 nsew power bidirectional
flabel metal4 s 98924 2128 99244 60432 0 FreeSans 1920 90 0 0 vccd1
port 43 nsew power bidirectional
flabel metal4 s 4868 59650 5188 101776 0 FreeSans 1920 90 0 0 vssd1
port 44 nsew ground bidirectional
flabel metal4 s 35588 59650 35908 101776 0 FreeSans 1920 90 0 0 vssd1
port 44 nsew ground bidirectional
flabel metal4 s 66308 59650 66628 101776 0 FreeSans 1920 90 0 0 vssd1
port 44 nsew ground bidirectional
flabel metal4 s 97028 59650 97348 101776 0 FreeSans 1920 90 0 0 vssd1
port 44 nsew ground bidirectional
flabel metal5 s 1056 6006 100880 6326 0 FreeSans 2560 0 0 0 vssd1
port 44 nsew ground bidirectional
flabel metal5 s 1056 36642 100880 36962 0 FreeSans 2560 0 0 0 vssd1
port 44 nsew ground bidirectional
flabel metal5 s 1056 67278 100880 67598 0 FreeSans 2560 0 0 0 vssd1
port 44 nsew ground bidirectional
flabel metal5 s 1056 97914 100880 98234 0 FreeSans 2560 0 0 0 vssd1
port 44 nsew ground bidirectional
flabel metal4 s 1668 2128 1828 60432 0 FreeSans 960 90 0 0 vssd1
port 44 nsew ground bidirectional
flabel metal4 s 99660 2128 99980 60432 0 FreeSans 1920 90 0 0 vssd1
port 44 nsew ground bidirectional
rlabel via4 95806 36142 95806 36142 0 vccd1
rlabel via4 95110 36802 95110 36802 0 vssd1
rlabel metal1 85836 60282 85836 60282 0 _000_
rlabel metal1 87676 60282 87676 60282 0 _001_
rlabel metal2 98486 40868 98486 40868 0 _002_
rlabel metal1 99820 29002 99820 29002 0 _003_
rlabel metal1 99636 27574 99636 27574 0 _004_
rlabel metal1 99130 23834 99130 23834 0 _005_
rlabel metal2 99406 23732 99406 23732 0 _006_
rlabel metal2 98854 19040 98854 19040 0 _007_
rlabel metal2 53222 76024 53222 76024 0 _008_
rlabel metal1 54142 74970 54142 74970 0 _009_
rlabel metal2 56902 76160 56902 76160 0 _010_
rlabel metal1 57914 74970 57914 74970 0 _011_
rlabel metal1 59984 74970 59984 74970 0 _012_
rlabel metal1 77464 60622 77464 60622 0 _013_
rlabel metal1 79120 60622 79120 60622 0 _014_
rlabel metal1 79488 60690 79488 60690 0 _015_
rlabel metal1 82011 60758 82011 60758 0 _016_
rlabel metal1 82340 60282 82340 60282 0 _017_
rlabel metal2 84042 60894 84042 60894 0 _018_
rlabel metal1 86013 60758 86013 60758 0 _019_
rlabel metal2 98394 42126 98394 42126 0 _020_
rlabel metal1 98578 35462 98578 35462 0 _021_
rlabel metal2 98394 32572 98394 32572 0 _022_
rlabel metal1 98670 25296 98670 25296 0 _023_
rlabel metal1 98709 24786 98709 24786 0 _024_
rlabel metal2 98486 21896 98486 21896 0 _025_
rlabel metal1 23283 61098 23283 61098 0 _026_
rlabel metal1 24242 60792 24242 60792 0 _027_
rlabel metal1 46138 74970 46138 74970 0 _028_
rlabel metal2 48254 76024 48254 76024 0 _029_
rlabel metal2 50002 76160 50002 76160 0 _030_
rlabel metal1 51520 74970 51520 74970 0 _031_
rlabel metal1 99809 26010 99809 26010 0 _032_
rlabel metal1 98532 40494 98532 40494 0 _033_
rlabel metal1 99636 27506 99636 27506 0 _034_
rlabel metal2 98302 24684 98302 24684 0 _035_
rlabel metal1 98716 22746 98716 22746 0 _036_
rlabel metal2 98670 20026 98670 20026 0 _037_
rlabel metal1 99498 22576 99498 22576 0 _038_
rlabel metal4 17470 3738 17470 3738 0 addr0[0]
rlabel metal4 18638 3874 18638 3874 0 addr0[1]
rlabel metal3 3703 27933 3703 27933 0 addr0[2]
rlabel metal3 1119 29308 1119 29308 0 addr0[3]
rlabel metal3 3703 30696 3703 30696 0 addr0[4]
rlabel metal3 3703 32396 3703 32396 0 addr0[5]
rlabel metal3 3059 33524 3059 33524 0 addr0[6]
rlabel metal3 3703 35224 3703 35224 0 addr0[7]
rlabel metal2 57086 59330 57086 59330 0 clk
rlabel metal1 55499 59942 55499 59942 0 clknet_0_clk
rlabel metal2 22402 59942 22402 59942 0 clknet_1_0__leaf_clk
rlabel metal2 77050 60656 77050 60656 0 clknet_1_1__leaf_clk
rlabel metal3 3703 9453 3703 9453 0 csb0
rlabel metal4 19806 3738 19806 3738 0 din0[0]
rlabel metal4 31486 3874 31486 3874 0 din0[10]
rlabel metal2 32890 1775 32890 1775 0 din0[11]
rlabel metal4 33822 3738 33822 3738 0 din0[12]
rlabel metal4 34990 3738 34990 3738 0 din0[13]
rlabel metal2 36110 1775 36110 1775 0 din0[14]
rlabel metal4 37326 3874 37326 3874 0 din0[15]
rlabel metal4 20974 3738 20974 3738 0 din0[1]
rlabel metal4 22142 3738 22142 3738 0 din0[2]
rlabel metal4 23310 3874 23310 3874 0 din0[3]
rlabel metal4 24478 3738 24478 3738 0 din0[4]
rlabel metal4 25646 3738 25646 3738 0 din0[5]
rlabel metal4 26814 3738 26814 3738 0 din0[6]
rlabel metal2 27738 2115 27738 2115 0 din0[7]
rlabel metal4 29164 3398 29164 3398 0 din0[8]
rlabel metal4 30318 3738 30318 3738 0 din0[9]
rlabel metal1 99636 26350 99636 26350 0 net1
rlabel metal2 43562 89556 43562 89556 0 net10
rlabel metal1 45448 101422 45448 101422 0 net11
rlabel metal1 47656 101422 47656 101422 0 net12
rlabel metal2 49726 89556 49726 89556 0 net13
rlabel metal1 51244 101422 51244 101422 0 net14
rlabel metal1 53176 101422 53176 101422 0 net15
rlabel metal1 55338 101422 55338 101422 0 net16
rlabel metal1 57408 101422 57408 101422 0 net17
rlabel metal1 57730 74834 57730 74834 0 net18
rlabel metal2 79258 60384 79258 60384 0 net19
rlabel metal2 21114 61574 21114 61574 0 net2
rlabel metal1 60490 74800 60490 74800 0 net20
rlabel metal3 96247 53738 96247 53738 0 net21
rlabel metal2 98486 18700 98486 18700 0 net22
rlabel metal1 85836 60078 85836 60078 0 net23
rlabel metal1 99682 29138 99682 29138 0 net24
rlabel metal1 87814 60146 87814 60146 0 net25
rlabel metal1 99406 27438 99406 27438 0 net26
rlabel metal1 59110 101422 59110 101422 0 net3
rlabel metal1 79718 61030 79718 61030 0 net4
rlabel metal2 96922 61744 96922 61744 0 net5
rlabel metal1 100234 60146 100234 60146 0 net6
rlabel metal2 100234 61030 100234 61030 0 net7
rlabel metal2 83858 60928 83858 60928 0 net8
rlabel metal2 1886 61302 1886 61302 0 net9
rlabel metal3 100886 25908 100886 25908 0 rst
rlabel metal3 751 61268 751 61268 0 sine_out[0]
rlabel metal2 58834 102527 58834 102527 0 sine_out[10]
rlabel via2 100418 62645 100418 62645 0 sine_out[11]
rlabel metal2 100418 62033 100418 62033 0 sine_out[12]
rlabel via2 100418 59925 100418 59925 0 sine_out[13]
rlabel metal2 100418 61421 100418 61421 0 sine_out[14]
rlabel via2 100418 60571 100418 60571 0 sine_out[15]
rlabel metal3 1096 61948 1096 61948 0 sine_out[1]
rlabel metal2 43378 102527 43378 102527 0 sine_out[2]
rlabel metal2 45310 102527 45310 102527 0 sine_out[3]
rlabel metal2 47978 102527 47978 102527 0 sine_out[4]
rlabel metal1 49726 101626 49726 101626 0 sine_out[5]
rlabel metal1 51060 101626 51060 101626 0 sine_out[6]
rlabel metal2 53038 102527 53038 102527 0 sine_out[7]
rlabel metal2 55706 102527 55706 102527 0 sine_out[8]
rlabel metal2 57638 102527 57638 102527 0 sine_out[9]
rlabel metal2 28198 59551 28198 59551 0 sine_out_temp\[0\]
rlabel metal1 57638 77418 57638 77418 0 sine_out_temp\[10\]
rlabel metal4 57563 57923 57563 57923 0 sine_out_temp\[11\]
rlabel metal4 60076 58127 60076 58127 0 sine_out_temp\[12\]
rlabel metal4 62652 58412 62652 58412 0 sine_out_temp\[13\]
rlabel metal4 65051 57787 65051 57787 0 sine_out_temp\[14\]
rlabel metal1 79534 61370 79534 61370 0 sine_out_temp\[15\]
rlabel metal2 24058 60452 24058 60452 0 sine_out_temp\[1\]
rlabel metal1 41768 77350 41768 77350 0 sine_out_temp\[2\]
rlabel metal4 37595 57923 37595 57923 0 sine_out_temp\[3\]
rlabel metal4 40158 58140 40158 58140 0 sine_out_temp\[4\]
rlabel metal4 42596 66831 42596 66831 0 sine_out_temp\[5\]
rlabel metal4 45083 57923 45083 57923 0 sine_out_temp\[6\]
rlabel metal1 51336 76806 51336 76806 0 sine_out_temp\[7\]
rlabel metal4 50075 57923 50075 57923 0 sine_out_temp\[8\]
rlabel metal2 55614 75701 55614 75701 0 sine_out_temp\[9\]
rlabel metal1 98348 44778 98348 44778 0 tcout\[0\]
rlabel metal1 98394 45050 98394 45050 0 tcout\[1\]
rlabel metal3 97405 19108 97405 19108 0 tcout\[2\]
rlabel metal1 98256 22678 98256 22678 0 tcout\[3\]
rlabel metal1 98532 22406 98532 22406 0 tcout\[4\]
rlabel metal1 97942 22746 97942 22746 0 tcout\[5\]
rlabel metal1 97934 21930 97934 21930 0 tcout\[6\]
rlabel metal1 98716 19278 98716 19278 0 tcout\[7\]
<< properties >>
string FIXED_BBOX 0 0 101962 104106
<< end >>
