module counter (clk,
    csb00,
    csb01,
    rst,
    addr00,
    addr01,
    din00,
    din01,
    sine_out);
 input clk;
 input csb00;
 input csb01;
 input rst;
 input [7:0] addr00;
 input [7:0] addr01;
 input [15:0] din00;
 input [15:0] din01;
 output [15:0] sine_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire net90;
 wire clknet_0_clk;
 wire \sine_out_temp0[0] ;
 wire \sine_out_temp0[10] ;
 wire \sine_out_temp0[11] ;
 wire \sine_out_temp0[12] ;
 wire \sine_out_temp0[13] ;
 wire \sine_out_temp0[14] ;
 wire \sine_out_temp0[15] ;
 wire \sine_out_temp0[1] ;
 wire \sine_out_temp0[2] ;
 wire \sine_out_temp0[3] ;
 wire \sine_out_temp0[4] ;
 wire \sine_out_temp0[5] ;
 wire \sine_out_temp0[6] ;
 wire \sine_out_temp0[7] ;
 wire \sine_out_temp0[8] ;
 wire \sine_out_temp0[9] ;
 wire \sine_out_temp1[0] ;
 wire \sine_out_temp1[10] ;
 wire \sine_out_temp1[11] ;
 wire \sine_out_temp1[12] ;
 wire \sine_out_temp1[13] ;
 wire \sine_out_temp1[14] ;
 wire \sine_out_temp1[15] ;
 wire \sine_out_temp1[1] ;
 wire \sine_out_temp1[2] ;
 wire \sine_out_temp1[3] ;
 wire \sine_out_temp1[4] ;
 wire \sine_out_temp1[5] ;
 wire \sine_out_temp1[6] ;
 wire \sine_out_temp1[7] ;
 wire \sine_out_temp1[8] ;
 wire \sine_out_temp1[9] ;
 wire \tcout[0] ;
 wire \tcout[1] ;
 wire \tcout[2] ;
 wire \tcout[3] ;
 wire \tcout[4] ;
 wire \tcout[5] ;
 wire \tcout[6] ;
 wire \tcout[7] ;
 wire \tcout[8] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;

 sky130_fd_sc_hd__inv_2 _061_ (.A(\tcout[0] ),
    .Y(_016_));
 sky130_fd_sc_hd__inv_2 _062_ (.A(net86),
    .Y(_025_));
 sky130_fd_sc_hd__mux2_1 _063_ (.A0(\sine_out_temp0[0] ),
    .A1(net83),
    .S(net84),
    .X(_000_));
 sky130_fd_sc_hd__mux2_1 _064_ (.A0(\sine_out_temp0[1] ),
    .A1(net76),
    .S(net84),
    .X(_007_));
 sky130_fd_sc_hd__mux2_1 _065_ (.A0(\sine_out_temp0[2] ),
    .A1(net75),
    .S(net84),
    .X(_008_));
 sky130_fd_sc_hd__mux2_1 _066_ (.A0(\sine_out_temp0[3] ),
    .A1(net74),
    .S(net84),
    .X(_009_));
 sky130_fd_sc_hd__mux2_1 _067_ (.A0(\sine_out_temp0[4] ),
    .A1(net73),
    .S(net84),
    .X(_010_));
 sky130_fd_sc_hd__mux2_1 _068_ (.A0(\sine_out_temp0[5] ),
    .A1(net72),
    .S(net84),
    .X(_011_));
 sky130_fd_sc_hd__mux2_1 _069_ (.A0(\sine_out_temp0[6] ),
    .A1(net71),
    .S(net84),
    .X(_012_));
 sky130_fd_sc_hd__mux2_1 _070_ (.A0(\sine_out_temp0[7] ),
    .A1(net70),
    .S(net84),
    .X(_013_));
 sky130_fd_sc_hd__mux2_1 _071_ (.A0(\sine_out_temp0[8] ),
    .A1(net69),
    .S(net84),
    .X(_014_));
 sky130_fd_sc_hd__mux2_1 _072_ (.A0(\sine_out_temp0[9] ),
    .A1(net68),
    .S(net84),
    .X(_015_));
 sky130_fd_sc_hd__mux2_1 _073_ (.A0(\sine_out_temp0[10] ),
    .A1(net82),
    .S(net85),
    .X(_001_));
 sky130_fd_sc_hd__mux2_1 _074_ (.A0(\sine_out_temp0[11] ),
    .A1(net81),
    .S(net85),
    .X(_002_));
 sky130_fd_sc_hd__mux2_1 _075_ (.A0(\sine_out_temp0[12] ),
    .A1(net80),
    .S(net85),
    .X(_003_));
 sky130_fd_sc_hd__mux2_1 _076_ (.A0(\sine_out_temp0[13] ),
    .A1(net79),
    .S(net85),
    .X(_004_));
 sky130_fd_sc_hd__mux2_1 _077_ (.A0(\sine_out_temp0[14] ),
    .A1(net78),
    .S(net85),
    .X(_005_));
 sky130_fd_sc_hd__mux2_1 _078_ (.A0(\sine_out_temp0[15] ),
    .A1(net77),
    .S(net85),
    .X(_006_));
 sky130_fd_sc_hd__xor2_1 _079_ (.A(\tcout[0] ),
    .B(\tcout[1] ),
    .X(_017_));
 sky130_fd_sc_hd__and3_1 _080_ (.A(\tcout[0] ),
    .B(\tcout[1] ),
    .C(\tcout[2] ),
    .X(_050_));
 sky130_fd_sc_hd__a21oi_1 _081_ (.A1(\tcout[0] ),
    .A2(\tcout[1] ),
    .B1(\tcout[2] ),
    .Y(_051_));
 sky130_fd_sc_hd__nor2_1 _082_ (.A(_050_),
    .B(_051_),
    .Y(_018_));
 sky130_fd_sc_hd__and4_2 _083_ (.A(\tcout[0] ),
    .B(\tcout[1] ),
    .C(\tcout[2] ),
    .D(\tcout[3] ),
    .X(_052_));
 sky130_fd_sc_hd__nor2_1 _084_ (.A(\tcout[3] ),
    .B(_050_),
    .Y(_053_));
 sky130_fd_sc_hd__nor2_1 _085_ (.A(_052_),
    .B(_053_),
    .Y(_019_));
 sky130_fd_sc_hd__xor2_1 _086_ (.A(\tcout[4] ),
    .B(_052_),
    .X(_020_));
 sky130_fd_sc_hd__and3_1 _087_ (.A(\tcout[4] ),
    .B(\tcout[5] ),
    .C(_052_),
    .X(_054_));
 sky130_fd_sc_hd__a21oi_1 _088_ (.A1(\tcout[4] ),
    .A2(_052_),
    .B1(\tcout[5] ),
    .Y(_055_));
 sky130_fd_sc_hd__nor2_1 _089_ (.A(_054_),
    .B(_055_),
    .Y(_021_));
 sky130_fd_sc_hd__xor2_1 _090_ (.A(\tcout[6] ),
    .B(_054_),
    .X(_022_));
 sky130_fd_sc_hd__and2_1 _091_ (.A(\tcout[6] ),
    .B(\tcout[7] ),
    .X(_056_));
 sky130_fd_sc_hd__and4_2 _092_ (.A(\tcout[4] ),
    .B(\tcout[5] ),
    .C(_052_),
    .D(_056_),
    .X(_057_));
 sky130_fd_sc_hd__a41o_1 _093_ (.A1(\tcout[4] ),
    .A2(\tcout[5] ),
    .A3(\tcout[6] ),
    .A4(_052_),
    .B1(\tcout[7] ),
    .X(_058_));
 sky130_fd_sc_hd__and2b_1 _094_ (.A_N(_057_),
    .B(_058_),
    .X(_023_));
 sky130_fd_sc_hd__xor2_1 _095_ (.A(net85),
    .B(_057_),
    .X(_024_));
 sky130_fd_sc_hd__inv_2 _096_ (.A(net87),
    .Y(_026_));
 sky130_fd_sc_hd__inv_2 _097_ (.A(net86),
    .Y(_027_));
 sky130_fd_sc_hd__inv_2 _098_ (.A(net86),
    .Y(_028_));
 sky130_fd_sc_hd__inv_2 _099_ (.A(net86),
    .Y(_029_));
 sky130_fd_sc_hd__inv_2 _100_ (.A(net86),
    .Y(_030_));
 sky130_fd_sc_hd__inv_2 _101_ (.A(net86),
    .Y(_031_));
 sky130_fd_sc_hd__inv_2 _102_ (.A(net87),
    .Y(_032_));
 sky130_fd_sc_hd__inv_2 _103_ (.A(net86),
    .Y(_033_));
 sky130_fd_sc_hd__inv_2 _104_ (.A(net87),
    .Y(_034_));
 sky130_fd_sc_hd__inv_2 _105_ (.A(net86),
    .Y(_035_));
 sky130_fd_sc_hd__inv_2 _106_ (.A(net87),
    .Y(_036_));
 sky130_fd_sc_hd__inv_2 _107_ (.A(net86),
    .Y(_037_));
 sky130_fd_sc_hd__inv_2 _108_ (.A(net87),
    .Y(_038_));
 sky130_fd_sc_hd__inv_2 _109_ (.A(net87),
    .Y(_039_));
 sky130_fd_sc_hd__inv_2 _110_ (.A(net86),
    .Y(_040_));
 sky130_fd_sc_hd__inv_2 _111_ (.A(net88),
    .Y(_041_));
 sky130_fd_sc_hd__inv_2 _112_ (.A(net88),
    .Y(_042_));
 sky130_fd_sc_hd__inv_2 _113_ (.A(net88),
    .Y(_043_));
 sky130_fd_sc_hd__inv_2 _114_ (.A(net88),
    .Y(_044_));
 sky130_fd_sc_hd__inv_2 _115_ (.A(net88),
    .Y(_045_));
 sky130_fd_sc_hd__inv_2 _116_ (.A(net88),
    .Y(_046_));
 sky130_fd_sc_hd__inv_2 _117_ (.A(net88),
    .Y(_047_));
 sky130_fd_sc_hd__inv_2 _118_ (.A(net88),
    .Y(_048_));
 sky130_fd_sc_hd__inv_2 _119_ (.A(net88),
    .Y(_049_));
 sky130_fd_sc_hd__dfrtp_1 _120_ (.CLK(clknet_2_2__leaf_clk),
    .D(_014_),
    .RESET_B(_025_),
    .Q(net66));
 sky130_fd_sc_hd__dfrtp_1 _121_ (.CLK(clknet_2_0__leaf_clk),
    .D(_015_),
    .RESET_B(_026_),
    .Q(net67));
 sky130_fd_sc_hd__dfrtp_1 _122_ (.CLK(clknet_2_1__leaf_clk),
    .D(_001_),
    .RESET_B(_027_),
    .Q(net53));
 sky130_fd_sc_hd__dfrtp_1 _123_ (.CLK(clknet_2_0__leaf_clk),
    .D(_002_),
    .RESET_B(_028_),
    .Q(net54));
 sky130_fd_sc_hd__dfrtp_1 _124_ (.CLK(clknet_2_1__leaf_clk),
    .D(_003_),
    .RESET_B(_029_),
    .Q(net55));
 sky130_fd_sc_hd__dfrtp_1 _125_ (.CLK(clknet_2_1__leaf_clk),
    .D(_004_),
    .RESET_B(_030_),
    .Q(net56));
 sky130_fd_sc_hd__dfrtp_1 _126_ (.CLK(clknet_2_3__leaf_clk),
    .D(_005_),
    .RESET_B(_031_),
    .Q(net57));
 sky130_fd_sc_hd__dfrtp_1 _127_ (.CLK(clknet_2_1__leaf_clk),
    .D(_006_),
    .RESET_B(_032_),
    .Q(net58));
 sky130_fd_sc_hd__dfrtp_4 _128_ (.CLK(clknet_2_3__leaf_clk),
    .D(_016_),
    .RESET_B(_033_),
    .Q(\tcout[0] ));
 sky130_fd_sc_hd__dfrtp_4 _129_ (.CLK(clknet_2_3__leaf_clk),
    .D(_017_),
    .RESET_B(_034_),
    .Q(\tcout[1] ));
 sky130_fd_sc_hd__dfrtp_4 _130_ (.CLK(clknet_2_1__leaf_clk),
    .D(_018_),
    .RESET_B(_035_),
    .Q(\tcout[2] ));
 sky130_fd_sc_hd__dfrtp_4 _131_ (.CLK(clknet_2_1__leaf_clk),
    .D(_019_),
    .RESET_B(_036_),
    .Q(\tcout[3] ));
 sky130_fd_sc_hd__dfrtp_4 _132_ (.CLK(clknet_2_1__leaf_clk),
    .D(_020_),
    .RESET_B(_037_),
    .Q(\tcout[4] ));
 sky130_fd_sc_hd__dfrtp_4 _133_ (.CLK(clknet_2_3__leaf_clk),
    .D(_021_),
    .RESET_B(_038_),
    .Q(\tcout[5] ));
 sky130_fd_sc_hd__dfrtp_4 _134_ (.CLK(clknet_2_1__leaf_clk),
    .D(_022_),
    .RESET_B(_039_),
    .Q(\tcout[6] ));
 sky130_fd_sc_hd__dfrtp_4 _135_ (.CLK(clknet_2_1__leaf_clk),
    .D(_023_),
    .RESET_B(_040_),
    .Q(\tcout[7] ));
 sky130_fd_sc_hd__dfrtp_1 _136_ (.CLK(clknet_2_2__leaf_clk),
    .D(_024_),
    .RESET_B(_041_),
    .Q(\tcout[8] ));
 sky130_fd_sc_hd__dfrtp_1 _137_ (.CLK(clknet_2_2__leaf_clk),
    .D(_000_),
    .RESET_B(_042_),
    .Q(net52));
 sky130_fd_sc_hd__dfrtp_1 _138_ (.CLK(clknet_2_0__leaf_clk),
    .D(_007_),
    .RESET_B(_043_),
    .Q(net59));
 sky130_fd_sc_hd__dfrtp_1 _139_ (.CLK(clknet_2_2__leaf_clk),
    .D(_008_),
    .RESET_B(_044_),
    .Q(net60));
 sky130_fd_sc_hd__dfrtp_1 _140_ (.CLK(clknet_2_0__leaf_clk),
    .D(_009_),
    .RESET_B(_045_),
    .Q(net61));
 sky130_fd_sc_hd__dfrtp_1 _141_ (.CLK(clknet_2_0__leaf_clk),
    .D(_010_),
    .RESET_B(_046_),
    .Q(net62));
 sky130_fd_sc_hd__dfrtp_1 _142_ (.CLK(clknet_2_0__leaf_clk),
    .D(_011_),
    .RESET_B(_047_),
    .Q(net63));
 sky130_fd_sc_hd__dfrtp_1 _143_ (.CLK(clknet_2_0__leaf_clk),
    .D(_012_),
    .RESET_B(_048_),
    .Q(net64));
 sky130_fd_sc_hd__dfrtp_1 _144_ (.CLK(clknet_2_3__leaf_clk),
    .D(_013_),
    .RESET_B(_049_),
    .Q(net65));
 sky130_fd_sc_hd__conb_1 mem_i1_90 (.LO(net90));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 ram256x16 mem_i0 (.csb0(net17),
    .csb1(net89),
    .clk0(clknet_2_0__leaf_clk),
    .clk1(clknet_2_1__leaf_clk),
    .addr0({net8,
    net7,
    net6,
    net5,
    net4,
    net3,
    net2,
    net1}),
    .addr1({\tcout[7] ,
    \tcout[6] ,
    \tcout[5] ,
    \tcout[4] ,
    \tcout[3] ,
    \tcout[2] ,
    \tcout[1] ,
    \tcout[0] }),
    .din0({net25,
    net24,
    net23,
    net22,
    net21,
    net20,
    net34,
    net33,
    net32,
    net31,
    net30,
    net29,
    net28,
    net27,
    net26,
    net19}),
    .dout1({\sine_out_temp0[15] ,
    \sine_out_temp0[14] ,
    \sine_out_temp0[13] ,
    \sine_out_temp0[12] ,
    \sine_out_temp0[11] ,
    \sine_out_temp0[10] ,
    \sine_out_temp0[9] ,
    \sine_out_temp0[8] ,
    \sine_out_temp0[7] ,
    \sine_out_temp0[6] ,
    \sine_out_temp0[5] ,
    \sine_out_temp0[4] ,
    \sine_out_temp0[3] ,
    \sine_out_temp0[2] ,
    \sine_out_temp0[1] ,
    \sine_out_temp0[0] }));
 ram256x16 mem_i1 (.csb0(net18),
    .csb1(net90),
    .clk0(clknet_2_2__leaf_clk),
    .clk1(clknet_2_3__leaf_clk),
    .addr0({net16,
    net15,
    net14,
    net13,
    net12,
    net11,
    net10,
    net9}),
    .addr1({\tcout[7] ,
    \tcout[6] ,
    \tcout[5] ,
    \tcout[4] ,
    \tcout[3] ,
    \tcout[2] ,
    \tcout[1] ,
    \tcout[0] }),
    .din0({net41,
    net40,
    net39,
    net38,
    net37,
    net36,
    net50,
    net49,
    net48,
    net47,
    net46,
    net45,
    net44,
    net43,
    net42,
    net35}),
    .dout1({\sine_out_temp1[15] ,
    \sine_out_temp1[14] ,
    \sine_out_temp1[13] ,
    \sine_out_temp1[12] ,
    \sine_out_temp1[11] ,
    \sine_out_temp1[10] ,
    \sine_out_temp1[9] ,
    \sine_out_temp1[8] ,
    \sine_out_temp1[7] ,
    \sine_out_temp1[6] ,
    \sine_out_temp1[5] ,
    \sine_out_temp1[4] ,
    \sine_out_temp1[3] ,
    \sine_out_temp1[2] ,
    \sine_out_temp1[1] ,
    \sine_out_temp1[0] }));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_117_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_118_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_119_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_120_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_228_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_229_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_2_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_2_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_2_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_2_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_2_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_2_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_2_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_2_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_2_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_2_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_2_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_2_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_2_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_2_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_2_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_2_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_2_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_2_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_2_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_2_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_2_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_2_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_2_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_2_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_2_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_2_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_2_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_2_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_2_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_2_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_2_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_2_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_2_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_2_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_2_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_2_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_2_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_2_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_2_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_2_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_2_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_2_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_2_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_2_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_2_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_2_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_2_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_2_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_2_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_2_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_2_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_2_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_2_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_2_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_2_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_2_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_2_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_2_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_2_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_2_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_2_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_2_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_2_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_2_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_2_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_2_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_2_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_2_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_2_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_2_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_2_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_2_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_2_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_2_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_2_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_2_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_2_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_2_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_2_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_2_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_2_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_2_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_2_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_2_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_2_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_2_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_2_Right_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_2_Right_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_2_Right_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_2_Right_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_2_Right_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_2_Right_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_2_Right_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_2_Right_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_2_Right_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_2_Right_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_2_Right_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_2_Right_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_2_Right_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_2_Right_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_2_Right_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_2_Right_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_2_Right_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_2_Right_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_2_Right_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_2_Right_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_2_Right_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_121_2_Right_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_122_2_Right_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_123_2_Right_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_124_2_Right_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_125_2_Right_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_126_2_Right_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_127_2_Right_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_128_2_Right_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_129_2_Right_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_130_2_Right_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_131_2_Right_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_132_2_Right_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_133_2_Right_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_134_2_Right_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_135_2_Right_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_136_2_Right_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_137_2_Right_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_138_2_Right_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_139_2_Right_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_140_2_Right_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_141_2_Right_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_142_2_Right_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_143_2_Right_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_144_2_Right_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_145_2_Right_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_146_2_Right_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_147_2_Right_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_148_2_Right_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_149_2_Right_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_150_2_Right_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_151_2_Right_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_152_2_Right_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_153_2_Right_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_154_2_Right_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_155_2_Right_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_156_2_Right_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_157_2_Right_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_158_2_Right_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_159_2_Right_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_160_2_Right_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_161_2_Right_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_162_2_Right_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_163_2_Right_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_164_2_Right_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_165_2_Right_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_166_2_Right_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_167_2_Right_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_168_2_Right_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_169_2_Right_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_170_2_Right_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_171_2_Right_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_172_2_Right_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_173_2_Right_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_174_2_Right_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_175_2_Right_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_176_2_Right_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_177_2_Right_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_178_2_Right_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_179_2_Right_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_180_2_Right_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_181_2_Right_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_182_2_Right_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_183_2_Right_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_184_2_Right_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_185_2_Right_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_186_2_Right_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_187_2_Right_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_188_2_Right_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_189_2_Right_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_190_2_Right_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_191_2_Right_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_192_2_Right_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_193_2_Right_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_194_2_Right_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_195_2_Right_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_196_2_Right_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_197_2_Right_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_198_2_Right_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_199_2_Right_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_200_2_Right_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_201_2_Right_203 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_202_2_Right_204 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_203_2_Right_205 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_204_2_Right_206 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_205_2_Right_207 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_206_2_Right_208 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_207_2_Right_209 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_208_2_Right_210 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_209_2_Right_211 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_210_2_Right_212 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_211_2_Right_213 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_212_2_Right_214 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_213_2_Right_215 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_214_2_Right_216 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_215_2_Right_217 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_216_2_Right_218 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_217_2_Right_219 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_218_2_Right_220 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_219_2_Right_221 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_220_2_Right_222 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_221_2_Right_223 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_222_2_Right_224 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_223_2_Right_225 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_224_2_Right_226 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_225_2_Right_227 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_226_2_Right_228 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_227_2_Right_229 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_230 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_231 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_232 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_233 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_234 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_235 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_236 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_237 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_238 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_239 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_1_Left_240 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_1_Left_241 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_1_Left_242 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_1_Left_243 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_1_Left_244 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_1_Left_245 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_1_Left_246 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_1_Left_247 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_1_Left_248 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_1_Left_249 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_1_Left_250 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_1_Left_251 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_1_Left_252 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_1_Left_253 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_1_Left_254 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_1_Left_255 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_1_Left_256 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_1_Left_257 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_1_Left_258 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_1_Left_259 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_1_Left_260 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_1_Left_261 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_1_Left_262 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_1_Left_263 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_1_Left_264 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_1_Left_265 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_1_Left_266 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_1_Left_267 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_1_Left_268 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_1_Left_269 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_1_Left_270 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_1_Left_271 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_1_Left_272 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_1_Left_273 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_1_Left_274 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_1_Left_275 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_1_Left_276 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_1_Left_277 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_1_Left_278 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_1_Left_279 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_1_Left_280 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_1_Left_281 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_1_Left_282 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_1_Left_283 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_1_Left_284 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_1_Left_285 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_1_Left_286 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_1_Left_287 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_1_Left_288 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_1_Left_289 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_1_Left_290 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_1_Left_291 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_1_Left_292 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_1_Left_293 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_1_Left_294 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_1_Left_295 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_1_Left_296 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_1_Left_297 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_1_Left_298 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_1_Left_299 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_1_Left_300 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_1_Left_301 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_1_Left_302 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_1_Left_303 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_1_Left_304 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_1_Left_305 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_1_Left_306 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_1_Left_307 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_1_Left_308 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_1_Left_309 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_1_Left_310 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_1_Left_311 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_1_Left_312 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_1_Left_313 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_1_Left_314 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_1_Left_315 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_1_Left_316 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_1_Left_317 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_1_Left_318 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_1_Left_319 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_1_Left_320 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_1_Left_321 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_1_Left_322 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_1_Left_323 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_1_Left_324 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_1_Left_325 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_1_Left_326 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_1_Left_327 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_1_Left_328 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_1_Left_329 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_1_Left_330 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_1_Left_331 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_1_Left_332 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_1_Left_333 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_1_Left_334 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_1_Left_335 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_1_Left_336 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_1_Left_337 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_1_Left_338 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_1_Left_339 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_1_Left_340 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_1_Left_341 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_1_Left_342 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_1_Left_343 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_1_Left_344 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_1_Left_345 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_121_1_Left_346 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_117_Left_347 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_118_Left_348 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_119_Left_349 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_120_Left_350 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_122_1_Left_351 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_123_1_Left_352 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_124_1_Left_353 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_125_1_Left_354 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_126_1_Left_355 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_127_1_Left_356 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_128_1_Left_357 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_129_1_Left_358 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_130_1_Left_359 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_131_1_Left_360 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_132_1_Left_361 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_133_1_Left_362 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_134_1_Left_363 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_135_1_Left_364 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_136_1_Left_365 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_137_1_Left_366 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_138_1_Left_367 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_139_1_Left_368 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_140_1_Left_369 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_141_1_Left_370 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_142_1_Left_371 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_143_1_Left_372 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_144_1_Left_373 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_145_1_Left_374 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_146_1_Left_375 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_147_1_Left_376 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_148_1_Left_377 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_149_1_Left_378 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_150_1_Left_379 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_151_1_Left_380 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_152_1_Left_381 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_153_1_Left_382 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_154_1_Left_383 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_155_1_Left_384 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_156_1_Left_385 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_157_1_Left_386 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_158_1_Left_387 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_159_1_Left_388 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_160_1_Left_389 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_161_1_Left_390 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_162_1_Left_391 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_163_1_Left_392 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_164_1_Left_393 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_165_1_Left_394 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_166_1_Left_395 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_167_1_Left_396 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_168_1_Left_397 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_169_1_Left_398 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_170_1_Left_399 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_171_1_Left_400 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_172_1_Left_401 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_173_1_Left_402 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_174_1_Left_403 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_175_1_Left_404 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_176_1_Left_405 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_177_1_Left_406 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_178_1_Left_407 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_179_1_Left_408 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_180_1_Left_409 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_181_1_Left_410 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_182_1_Left_411 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_183_1_Left_412 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_184_1_Left_413 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_185_1_Left_414 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_186_1_Left_415 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_187_1_Left_416 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_188_1_Left_417 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_189_1_Left_418 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_190_1_Left_419 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_191_1_Left_420 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_192_1_Left_421 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_193_1_Left_422 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_194_1_Left_423 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_195_1_Left_424 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_196_1_Left_425 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_197_1_Left_426 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_198_1_Left_427 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_199_1_Left_428 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_200_1_Left_429 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_201_1_Left_430 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_202_1_Left_431 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_203_1_Left_432 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_204_1_Left_433 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_205_1_Left_434 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_206_1_Left_435 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_207_1_Left_436 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_208_1_Left_437 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_209_1_Left_438 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_210_1_Left_439 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_211_1_Left_440 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_212_1_Left_441 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_213_1_Left_442 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_214_1_Left_443 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_215_1_Left_444 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_216_1_Left_445 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_217_1_Left_446 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_218_1_Left_447 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_219_1_Left_448 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_220_1_Left_449 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_221_1_Left_450 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_222_1_Left_451 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_223_1_Left_452 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_224_1_Left_453 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_225_1_Left_454 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_226_1_Left_455 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_227_1_Left_456 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_228_Left_457 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_229_Left_458 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_1_Left_459 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_2_Left_460 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_2_Left_461 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_2_Left_462 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_2_Left_463 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_2_Left_464 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_2_Left_465 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_2_Left_466 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_2_Left_467 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_2_Left_468 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_2_Left_469 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_2_Left_470 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_2_Left_471 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_2_Left_472 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_2_Left_473 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_2_Left_474 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_2_Left_475 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_2_Left_476 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_2_Left_477 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_2_Left_478 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_2_Left_479 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_2_Left_480 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_2_Left_481 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_2_Left_482 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_2_Left_483 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_2_Left_484 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_2_Left_485 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_2_Left_486 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_2_Left_487 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_2_Left_488 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_2_Left_489 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_2_Left_490 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_2_Left_491 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_2_Left_492 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_2_Left_493 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_2_Left_494 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_2_Left_495 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_2_Left_496 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_2_Left_497 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_2_Left_498 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_2_Left_499 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_2_Left_500 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_2_Left_501 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_2_Left_502 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_2_Left_503 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_2_Left_504 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_2_Left_505 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_2_Left_506 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_2_Left_507 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_2_Left_508 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_2_Left_509 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_2_Left_510 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_2_Left_511 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_2_Left_512 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_2_Left_513 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_2_Left_514 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_2_Left_515 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_2_Left_516 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_2_Left_517 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_2_Left_518 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_2_Left_519 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_2_Left_520 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_2_Left_521 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_2_Left_522 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_2_Left_523 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_2_Left_524 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_2_Left_525 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_2_Left_526 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_2_Left_527 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_2_Left_528 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_2_Left_529 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_2_Left_530 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_2_Left_531 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_2_Left_532 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_2_Left_533 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_2_Left_534 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_2_Left_535 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_2_Left_536 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_2_Left_537 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_2_Left_538 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_2_Left_539 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_2_Left_540 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_2_Left_541 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_2_Left_542 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_2_Left_543 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_2_Left_544 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_2_Left_545 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_2_Left_546 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_2_Left_547 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_2_Left_548 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_2_Left_549 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_2_Left_550 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_2_Left_551 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_2_Left_552 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_2_Left_553 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_2_Left_554 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_2_Left_555 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_2_Left_556 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_2_Left_557 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_2_Left_558 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_2_Left_559 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_2_Left_560 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_2_Left_561 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_2_Left_562 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_2_Left_563 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_2_Left_564 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_2_Left_565 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_2_Left_566 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_1_Right_567 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_1_Right_568 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_1_Right_569 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_1_Right_570 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_1_Right_571 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_1_Right_572 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_1_Right_573 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_1_Right_574 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_1_Right_575 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_1_Right_576 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_1_Right_577 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_1_Right_578 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_1_Right_579 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_1_Right_580 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_1_Right_581 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_1_Right_582 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_1_Right_583 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_1_Right_584 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_1_Right_585 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_1_Right_586 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_1_Right_587 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_1_Right_588 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_1_Right_589 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_1_Right_590 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_1_Right_591 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_1_Right_592 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_1_Right_593 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_1_Right_594 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_1_Right_595 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_1_Right_596 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_1_Right_597 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_1_Right_598 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_1_Right_599 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_1_Right_600 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_1_Right_601 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_1_Right_602 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_1_Right_603 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_1_Right_604 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_1_Right_605 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_1_Right_606 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_1_Right_607 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_1_Right_608 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_1_Right_609 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_1_Right_610 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_1_Right_611 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_1_Right_612 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_1_Right_613 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_1_Right_614 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_1_Right_615 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_1_Right_616 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_1_Right_617 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_1_Right_618 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_1_Right_619 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_1_Right_620 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_1_Right_621 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_1_Right_622 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_1_Right_623 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_1_Right_624 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_1_Right_625 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_1_Right_626 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_1_Right_627 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_1_Right_628 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_1_Right_629 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_1_Right_630 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_1_Right_631 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_1_Right_632 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_1_Right_633 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_1_Right_634 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_1_Right_635 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_1_Right_636 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_1_Right_637 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_1_Right_638 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_1_Right_639 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_1_Right_640 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_1_Right_641 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_1_Right_642 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_1_Right_643 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_1_Right_644 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_1_Right_645 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_1_Right_646 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_1_Right_647 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_1_Right_648 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_1_Right_649 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_1_Right_650 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_1_Right_651 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_1_Right_652 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_1_Right_653 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_1_Right_654 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_1_Right_655 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_1_Right_656 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_1_Right_657 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_1_Right_658 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_1_Right_659 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_1_Right_660 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_1_Right_661 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_1_Right_662 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_1_Right_663 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_1_Right_664 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_1_Right_665 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_1_Right_666 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_1_Right_667 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_1_Right_668 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_1_Right_669 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_1_Right_670 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_1_Right_671 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_1_Right_672 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_1_Right_673 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_121_2_Left_674 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_122_2_Left_675 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_123_2_Left_676 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_124_2_Left_677 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_125_2_Left_678 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_126_2_Left_679 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_127_2_Left_680 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_128_2_Left_681 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_129_2_Left_682 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_130_2_Left_683 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_131_2_Left_684 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_132_2_Left_685 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_133_2_Left_686 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_134_2_Left_687 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_135_2_Left_688 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_136_2_Left_689 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_137_2_Left_690 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_138_2_Left_691 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_139_2_Left_692 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_140_2_Left_693 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_141_2_Left_694 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_142_2_Left_695 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_143_2_Left_696 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_144_2_Left_697 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_145_2_Left_698 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_146_2_Left_699 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_147_2_Left_700 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_148_2_Left_701 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_149_2_Left_702 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_150_2_Left_703 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_151_2_Left_704 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_152_2_Left_705 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_153_2_Left_706 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_154_2_Left_707 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_155_2_Left_708 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_156_2_Left_709 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_157_2_Left_710 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_158_2_Left_711 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_159_2_Left_712 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_160_2_Left_713 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_161_2_Left_714 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_162_2_Left_715 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_163_2_Left_716 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_164_2_Left_717 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_165_2_Left_718 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_166_2_Left_719 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_167_2_Left_720 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_168_2_Left_721 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_169_2_Left_722 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_170_2_Left_723 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_171_2_Left_724 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_172_2_Left_725 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_173_2_Left_726 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_174_2_Left_727 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_175_2_Left_728 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_176_2_Left_729 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_177_2_Left_730 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_178_2_Left_731 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_179_2_Left_732 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_180_2_Left_733 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_181_2_Left_734 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_182_2_Left_735 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_183_2_Left_736 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_184_2_Left_737 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_185_2_Left_738 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_186_2_Left_739 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_187_2_Left_740 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_188_2_Left_741 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_189_2_Left_742 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_190_2_Left_743 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_191_2_Left_744 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_192_2_Left_745 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_193_2_Left_746 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_194_2_Left_747 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_195_2_Left_748 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_196_2_Left_749 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_197_2_Left_750 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_198_2_Left_751 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_199_2_Left_752 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_200_2_Left_753 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_201_2_Left_754 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_202_2_Left_755 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_203_2_Left_756 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_204_2_Left_757 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_205_2_Left_758 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_206_2_Left_759 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_207_2_Left_760 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_208_2_Left_761 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_209_2_Left_762 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_210_2_Left_763 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_211_2_Left_764 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_212_2_Left_765 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_213_2_Left_766 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_214_2_Left_767 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_215_2_Left_768 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_216_2_Left_769 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_217_2_Left_770 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_218_2_Left_771 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_219_2_Left_772 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_220_2_Left_773 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_221_2_Left_774 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_222_2_Left_775 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_223_2_Left_776 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_224_2_Left_777 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_225_2_Left_778 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_226_2_Left_779 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_227_2_Left_780 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_121_1_Right_781 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_122_1_Right_782 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_123_1_Right_783 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_124_1_Right_784 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_125_1_Right_785 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_126_1_Right_786 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_127_1_Right_787 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_128_1_Right_788 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_129_1_Right_789 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_130_1_Right_790 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_131_1_Right_791 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_132_1_Right_792 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_133_1_Right_793 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_134_1_Right_794 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_135_1_Right_795 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_136_1_Right_796 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_137_1_Right_797 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_138_1_Right_798 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_139_1_Right_799 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_140_1_Right_800 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_141_1_Right_801 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_142_1_Right_802 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_143_1_Right_803 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_144_1_Right_804 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_145_1_Right_805 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_146_1_Right_806 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_147_1_Right_807 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_148_1_Right_808 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_149_1_Right_809 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_150_1_Right_810 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_151_1_Right_811 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_152_1_Right_812 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_153_1_Right_813 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_154_1_Right_814 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_155_1_Right_815 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_156_1_Right_816 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_157_1_Right_817 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_158_1_Right_818 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_159_1_Right_819 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_160_1_Right_820 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_161_1_Right_821 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_162_1_Right_822 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_163_1_Right_823 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_164_1_Right_824 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_165_1_Right_825 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_166_1_Right_826 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_167_1_Right_827 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_168_1_Right_828 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_169_1_Right_829 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_170_1_Right_830 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_171_1_Right_831 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_172_1_Right_832 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_173_1_Right_833 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_174_1_Right_834 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_175_1_Right_835 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_176_1_Right_836 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_177_1_Right_837 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_178_1_Right_838 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_179_1_Right_839 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_180_1_Right_840 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_181_1_Right_841 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_182_1_Right_842 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_183_1_Right_843 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_184_1_Right_844 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_185_1_Right_845 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_186_1_Right_846 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_187_1_Right_847 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_188_1_Right_848 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_189_1_Right_849 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_190_1_Right_850 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_191_1_Right_851 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_192_1_Right_852 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_193_1_Right_853 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_194_1_Right_854 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_195_1_Right_855 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_196_1_Right_856 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_197_1_Right_857 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_198_1_Right_858 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_199_1_Right_859 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_200_1_Right_860 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_201_1_Right_861 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_202_1_Right_862 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_203_1_Right_863 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_204_1_Right_864 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_205_1_Right_865 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_206_1_Right_866 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_207_1_Right_867 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_208_1_Right_868 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_209_1_Right_869 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_210_1_Right_870 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_211_1_Right_871 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_212_1_Right_872 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_213_1_Right_873 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_214_1_Right_874 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_215_1_Right_875 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_216_1_Right_876 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_217_1_Right_877 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_218_1_Right_878 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_219_1_Right_879 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_220_1_Right_880 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_221_1_Right_881 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_222_1_Right_882 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_223_1_Right_883 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_224_1_Right_884 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_225_1_Right_885 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_226_1_Right_886 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_227_1_Right_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_1_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_1_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_1_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_1_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_1_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_1_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_1_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_1_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_1_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_1_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_1_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_1_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_1_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_1_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_1_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_1_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_1_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_1_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_1_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_1_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_1_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_1_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_1_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_1_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_1_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_1_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_1_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_1_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_1_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_1_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_1_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_1_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_1_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_1_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_1_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_1_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_1_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_1_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_1_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_1_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_1_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_1_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_1_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_1_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_1_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_1_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_1_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_1_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_1_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_1_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_1_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_1_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_1_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_1_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_1_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_1_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_1_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_1_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_1_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_1_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_1_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_1_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_1_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_1_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_1_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_1_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_1_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_1_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_1_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_1_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_1_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_1_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_1_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_1_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_1_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_1_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_1_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_1_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_1_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_1_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_1_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_1_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_1_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_1_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_1_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_1_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_1_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_1_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_1_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_1_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_1_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_1_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_1_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_1_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_1_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_1_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_1_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_1_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_2_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_2_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_2_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_2_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_2_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_2_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_2_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_2_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_2_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_2_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_2_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_2_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_2_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_2_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_2_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_2_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_2_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_2_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_2_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_2_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_2_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_2_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_2_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_2_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_2_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_2_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_2_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_2_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_2_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_2_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_2_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_2_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_2_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_2_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_2_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_2_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_2_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_2_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_2_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_2_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_2_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_2_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_2_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_2_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_2_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_2_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_2_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_2_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_2_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_2_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_2_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_2_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_2_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_2_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_2_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_2_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_2_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_2_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_2_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_2_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_2_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_2_1659 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(addr00[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(addr00[1]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(addr00[2]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(addr00[3]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(addr00[4]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(addr00[5]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(addr00[6]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(addr00[7]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_2 input9 (.A(addr01[0]),
    .X(net9));
 sky130_fd_sc_hd__dlymetal6s2s_1 input10 (.A(addr01[1]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(addr01[2]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(addr01[3]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(addr01[4]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(addr01[5]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(addr01[6]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(addr01[7]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(csb00),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(csb01),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(din00[0]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(din00[10]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(din00[11]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(din00[12]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(din00[13]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(din00[14]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(din00[15]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(din00[1]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(din00[2]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(din00[3]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(din00[4]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(din00[5]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(din00[6]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(din00[7]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(din00[8]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(din00[9]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_2 input35 (.A(din01[0]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_2 input36 (.A(din01[10]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_2 input37 (.A(din01[11]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_2 input38 (.A(din01[12]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_2 input39 (.A(din01[13]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_2 input40 (.A(din01[14]),
    .X(net40));
 sky130_fd_sc_hd__buf_2 input41 (.A(din01[15]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_2 input42 (.A(din01[1]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_2 input43 (.A(din01[2]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_2 input44 (.A(din01[3]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_2 input45 (.A(din01[4]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_2 input46 (.A(din01[5]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_2 input47 (.A(din01[6]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_2 input48 (.A(din01[7]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_2 input49 (.A(din01[8]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_2 input50 (.A(din01[9]),
    .X(net50));
 sky130_fd_sc_hd__buf_1 input51 (.A(rst),
    .X(net51));
 sky130_fd_sc_hd__buf_2 output52 (.A(net52),
    .X(sine_out[0]));
 sky130_fd_sc_hd__buf_2 output53 (.A(net53),
    .X(sine_out[10]));
 sky130_fd_sc_hd__buf_2 output54 (.A(net54),
    .X(sine_out[11]));
 sky130_fd_sc_hd__buf_2 output55 (.A(net55),
    .X(sine_out[12]));
 sky130_fd_sc_hd__buf_2 output56 (.A(net56),
    .X(sine_out[13]));
 sky130_fd_sc_hd__buf_2 output57 (.A(net57),
    .X(sine_out[14]));
 sky130_fd_sc_hd__buf_2 output58 (.A(net58),
    .X(sine_out[15]));
 sky130_fd_sc_hd__buf_2 output59 (.A(net59),
    .X(sine_out[1]));
 sky130_fd_sc_hd__buf_2 output60 (.A(net60),
    .X(sine_out[2]));
 sky130_fd_sc_hd__buf_2 output61 (.A(net61),
    .X(sine_out[3]));
 sky130_fd_sc_hd__buf_2 output62 (.A(net62),
    .X(sine_out[4]));
 sky130_fd_sc_hd__buf_2 output63 (.A(net63),
    .X(sine_out[5]));
 sky130_fd_sc_hd__buf_2 output64 (.A(net64),
    .X(sine_out[6]));
 sky130_fd_sc_hd__buf_2 output65 (.A(net65),
    .X(sine_out[7]));
 sky130_fd_sc_hd__buf_2 output66 (.A(net66),
    .X(sine_out[8]));
 sky130_fd_sc_hd__buf_2 output67 (.A(net67),
    .X(sine_out[9]));
 sky130_fd_sc_hd__clkbuf_2 wire68 (.A(\sine_out_temp1[9] ),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_2 wire69 (.A(\sine_out_temp1[8] ),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_2 wire70 (.A(\sine_out_temp1[7] ),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_2 wire71 (.A(\sine_out_temp1[6] ),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_2 wire72 (.A(\sine_out_temp1[5] ),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_2 wire73 (.A(\sine_out_temp1[4] ),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_2 wire74 (.A(\sine_out_temp1[3] ),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_2 wire75 (.A(\sine_out_temp1[2] ),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_2 wire76 (.A(\sine_out_temp1[1] ),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_2 wire77 (.A(\sine_out_temp1[15] ),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_2 wire78 (.A(\sine_out_temp1[14] ),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_2 wire79 (.A(\sine_out_temp1[13] ),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_2 wire80 (.A(\sine_out_temp1[12] ),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_2 wire81 (.A(\sine_out_temp1[11] ),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_2 wire82 (.A(\sine_out_temp1[10] ),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_2 wire83 (.A(\sine_out_temp1[0] ),
    .X(net83));
 sky130_fd_sc_hd__buf_4 fanout84 (.A(\tcout[8] ),
    .X(net84));
 sky130_fd_sc_hd__buf_2 fanout85 (.A(\tcout[8] ),
    .X(net85));
 sky130_fd_sc_hd__buf_4 fanout86 (.A(net87),
    .X(net86));
 sky130_fd_sc_hd__buf_4 fanout87 (.A(net88),
    .X(net87));
 sky130_fd_sc_hd__buf_6 fanout88 (.A(net51),
    .X(net88));
 sky130_fd_sc_hd__conb_1 mem_i0_89 (.LO(net89));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload0 (.A(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload1 (.A(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__bufinv_16 clkload2 (.A(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__124__D (.DIODE(_003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__075__X (.DIODE(_003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__126__D (.DIODE(_005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__077__X (.DIODE(_005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__141__D (.DIODE(_010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__067__X (.DIODE(_010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__142__D (.DIODE(_011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__068__X (.DIODE(_011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__082__B (.DIODE(_051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__081__Y (.DIODE(_051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__093__A4 (.DIODE(_052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__092__C (.DIODE(_052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__088__A2 (.DIODE(_052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__087__C (.DIODE(_052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__086__B (.DIODE(_052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__085__A (.DIODE(_052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__083__X (.DIODE(_052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__095__B (.DIODE(_057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__094__A_N (.DIODE(_057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__092__X (.DIODE(_057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__094__B (.DIODE(_058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__093__X (.DIODE(_058_));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(addr00[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(addr00[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(addr00[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(addr00[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(addr00[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(addr00[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(addr00[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(addr00[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(addr01[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(addr01[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(addr01[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(addr01[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(addr01[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(addr01[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(addr01[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(addr01[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(csb00));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(csb01));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(din00[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(din00[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(din00[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(din00[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(din00[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(din00[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(din00[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(din00[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(din00[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(din00[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(din00[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(din00[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(din00[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(din00[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(din00[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(din00[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(din01[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(din01[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(din01[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(din01[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(din01[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(din01[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_A (.DIODE(din01[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_A (.DIODE(din01[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_A (.DIODE(din01[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_A (.DIODE(din01[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_A (.DIODE(din01[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_A (.DIODE(din01[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_A (.DIODE(din01[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_A (.DIODE(din01[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_A (.DIODE(din01[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_A (.DIODE(din01[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_A (.DIODE(rst));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_dout1[7]  (.DIODE(\sine_out_temp0[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__070__A0 (.DIODE(\sine_out_temp0[7] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_addr1[0]  (.DIODE(\tcout[0] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_addr1[0]  (.DIODE(\tcout[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__128__Q (.DIODE(\tcout[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__083__A (.DIODE(\tcout[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__081__A1 (.DIODE(\tcout[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__080__A (.DIODE(\tcout[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__079__A (.DIODE(\tcout[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__061__A (.DIODE(\tcout[0] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_addr1[1]  (.DIODE(\tcout[1] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_addr1[1]  (.DIODE(\tcout[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__129__Q (.DIODE(\tcout[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__083__B (.DIODE(\tcout[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__081__A2 (.DIODE(\tcout[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__080__B (.DIODE(\tcout[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__079__B (.DIODE(\tcout[1] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_addr1[2]  (.DIODE(\tcout[2] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_addr1[2]  (.DIODE(\tcout[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__130__Q (.DIODE(\tcout[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__083__C (.DIODE(\tcout[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__081__B1 (.DIODE(\tcout[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__080__C (.DIODE(\tcout[2] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_addr1[3]  (.DIODE(\tcout[3] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_addr1[3]  (.DIODE(\tcout[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__131__Q (.DIODE(\tcout[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__084__A (.DIODE(\tcout[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__083__D (.DIODE(\tcout[3] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_addr1[4]  (.DIODE(\tcout[4] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_addr1[4]  (.DIODE(\tcout[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__132__Q (.DIODE(\tcout[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__093__A1 (.DIODE(\tcout[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__092__A (.DIODE(\tcout[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__088__A1 (.DIODE(\tcout[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__087__A (.DIODE(\tcout[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__086__A (.DIODE(\tcout[4] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_addr1[5]  (.DIODE(\tcout[5] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_addr1[5]  (.DIODE(\tcout[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__133__Q (.DIODE(\tcout[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__093__A2 (.DIODE(\tcout[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__092__B (.DIODE(\tcout[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__088__B1 (.DIODE(\tcout[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__087__B (.DIODE(\tcout[5] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_addr1[6]  (.DIODE(\tcout[6] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_addr1[6]  (.DIODE(\tcout[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__134__Q (.DIODE(\tcout[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__093__A3 (.DIODE(\tcout[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__091__A (.DIODE(\tcout[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__090__A (.DIODE(\tcout[6] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_addr1[7]  (.DIODE(\tcout[7] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i0_addr1[7]  (.DIODE(\tcout[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__135__Q (.DIODE(\tcout[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__093__B1 (.DIODE(\tcout[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__091__B (.DIODE(\tcout[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_X (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_addr0[0]  (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_X (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_addr0[1]  (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_X (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_din0[0]  (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_X (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_din0[10]  (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_X (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_din0[11]  (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_X (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_din0[12]  (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_X (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_din0[13]  (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_X (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_din0[14]  (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_X (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_din0[15]  (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_X (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_din0[1]  (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_X (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_din0[2]  (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_X (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_din0[3]  (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_X (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_din0[4]  (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_X (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_din0[5]  (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_X (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_din0[6]  (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_X (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_din0[7]  (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_X (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_din0[8]  (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_X (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mem_i1_din0[9]  (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_output52_A (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__137__Q (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_output53_A (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__122__Q (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_output54_A (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__123__Q (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_output56_A (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__125__Q (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_output59_A (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__138__Q (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_output60_A (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__139__Q (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_output61_A (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__140__Q (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_output62_A (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__141__Q (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_output63_A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__142__Q (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_output64_A (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__143__Q (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_output65_A (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__144__Q (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_output66_A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__120__Q (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_output67_A (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__121__Q (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire68_X (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__072__A1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire69_X (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__071__A1 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire70_X (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__070__A1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire71_X (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__069__A1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire72_X (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__068__A1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire73_X (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__067__A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire74_X (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__066__A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire75_X (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__065__A1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire76_X (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__064__A1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire77_X (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__078__A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire78_X (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__077__A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire79_X (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__076__A1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire80_X (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__075__A1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire81_X (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__074__A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire82_X (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__073__A1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire83_X (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__063__A1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout84_X (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__072__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__071__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__070__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__069__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__068__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__067__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__066__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__065__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__064__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__063__S (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout87_X (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout86_A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__096__A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__104__A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__106__A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__109__A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__108__A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__102__A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout88_X (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__111__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__119__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout87_A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__118__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__117__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__116__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__115__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__114__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__113__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__112__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkload0_A (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__121__CLK (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__123__CLK (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__138__CLK (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__140__CLK (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__141__CLK (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__142__CLK (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__143__CLK (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_mem_i0_clk0 (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0__f_clk_X (.DIODE(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__122__CLK (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__124__CLK (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__125__CLK (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__127__CLK (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__130__CLK (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__131__CLK (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__132__CLK (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__134__CLK (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__135__CLK (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_mem_i0_clk1 (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f_clk_X (.DIODE(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkload1_A (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__120__CLK (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__136__CLK (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__137__CLK (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__139__CLK (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_mem_i1_clk0 (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f_clk_X (.DIODE(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkload2_A (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__126__CLK (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__128__CLK (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__129__CLK (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__133__CLK (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__144__CLK (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_mem_i1_clk1 (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f_clk_X (.DIODE(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_015_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(\sine_out_temp0[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(\sine_out_temp0[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(\sine_out_temp0[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(\sine_out_temp0[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(\sine_out_temp0[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(\sine_out_temp0[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(\sine_out_temp0[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(_007_));
endmodule
