module counter (clk,
    csb0,
    rst,
    addr0,
    din0,
    sine_out);
 input clk;
 input csb0;
 input rst;
 input [7:0] addr0;
 input [15:0] din0;
 output [15:0] sine_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire \sine_out_temp[0] ;
 wire \sine_out_temp[10] ;
 wire \sine_out_temp[11] ;
 wire \sine_out_temp[12] ;
 wire \sine_out_temp[13] ;
 wire \sine_out_temp[14] ;
 wire \sine_out_temp[15] ;
 wire \sine_out_temp[1] ;
 wire \sine_out_temp[2] ;
 wire \sine_out_temp[3] ;
 wire \sine_out_temp[4] ;
 wire \sine_out_temp[5] ;
 wire \sine_out_temp[6] ;
 wire \sine_out_temp[7] ;
 wire \sine_out_temp[8] ;
 wire \sine_out_temp[9] ;
 wire \tcout[0] ;
 wire \tcout[1] ;
 wire \tcout[2] ;
 wire \tcout[3] ;
 wire \tcout[4] ;
 wire \tcout[5] ;
 wire \tcout[6] ;
 wire \tcout[7] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;

 sky130_fd_sc_hd__inv_2 _040_ (.A(\tcout[0] ),
    .Y(_000_));
 sky130_fd_sc_hd__inv_2 _041_ (.A(net18),
    .Y(_008_));
 sky130_fd_sc_hd__xor2_1 _042_ (.A(\tcout[0] ),
    .B(\tcout[1] ),
    .X(_001_));
 sky130_fd_sc_hd__and3_2 _043_ (.A(\tcout[0] ),
    .B(\tcout[1] ),
    .C(\tcout[2] ),
    .X(_032_));
 sky130_fd_sc_hd__a21oi_1 _044_ (.A1(\tcout[0] ),
    .A2(\tcout[1] ),
    .B1(\tcout[2] ),
    .Y(_033_));
 sky130_fd_sc_hd__nor2_1 _045_ (.A(_032_),
    .B(_033_),
    .Y(_002_));
 sky130_fd_sc_hd__nand2_1 _046_ (.A(\tcout[3] ),
    .B(_032_),
    .Y(_034_));
 sky130_fd_sc_hd__xor2_1 _047_ (.A(\tcout[3] ),
    .B(_032_),
    .X(_003_));
 sky130_fd_sc_hd__and3_1 _048_ (.A(\tcout[3] ),
    .B(\tcout[4] ),
    .C(_032_),
    .X(_035_));
 sky130_fd_sc_hd__xnor2_1 _049_ (.A(\tcout[4] ),
    .B(_034_),
    .Y(_004_));
 sky130_fd_sc_hd__and3_1 _050_ (.A(\tcout[3] ),
    .B(\tcout[4] ),
    .C(\tcout[5] ),
    .X(_036_));
 sky130_fd_sc_hd__o2bb2a_1 _051_ (.A1_N(_032_),
    .A2_N(_036_),
    .B1(_035_),
    .B2(\tcout[5] ),
    .X(_005_));
 sky130_fd_sc_hd__and3_1 _052_ (.A(\tcout[6] ),
    .B(_032_),
    .C(_036_),
    .X(_037_));
 sky130_fd_sc_hd__a21oi_1 _053_ (.A1(_032_),
    .A2(_036_),
    .B1(\tcout[6] ),
    .Y(_038_));
 sky130_fd_sc_hd__nor2_1 _054_ (.A(_037_),
    .B(_038_),
    .Y(_006_));
 sky130_fd_sc_hd__xor2_1 _055_ (.A(\tcout[7] ),
    .B(_037_),
    .X(_007_));
 sky130_fd_sc_hd__inv_2 _056_ (.A(net18),
    .Y(_009_));
 sky130_fd_sc_hd__inv_2 _057_ (.A(net18),
    .Y(_010_));
 sky130_fd_sc_hd__inv_2 _058_ (.A(net18),
    .Y(_011_));
 sky130_fd_sc_hd__inv_2 _059_ (.A(net19),
    .Y(_012_));
 sky130_fd_sc_hd__inv_2 _060_ (.A(net19),
    .Y(_013_));
 sky130_fd_sc_hd__inv_2 _061_ (.A(net19),
    .Y(_014_));
 sky130_fd_sc_hd__inv_2 _062_ (.A(net19),
    .Y(_015_));
 sky130_fd_sc_hd__inv_2 _063_ (.A(net19),
    .Y(_016_));
 sky130_fd_sc_hd__inv_2 _064_ (.A(net19),
    .Y(_017_));
 sky130_fd_sc_hd__inv_2 _065_ (.A(net20),
    .Y(_018_));
 sky130_fd_sc_hd__inv_2 _066_ (.A(net20),
    .Y(_019_));
 sky130_fd_sc_hd__inv_2 _067_ (.A(net20),
    .Y(_020_));
 sky130_fd_sc_hd__inv_2 _068_ (.A(net20),
    .Y(_021_));
 sky130_fd_sc_hd__inv_2 _069_ (.A(net20),
    .Y(_022_));
 sky130_fd_sc_hd__inv_2 _070_ (.A(net20),
    .Y(_023_));
 sky130_fd_sc_hd__inv_2 _071_ (.A(net20),
    .Y(_024_));
 sky130_fd_sc_hd__inv_2 _072_ (.A(net20),
    .Y(_025_));
 sky130_fd_sc_hd__inv_2 _073_ (.A(net18),
    .Y(_026_));
 sky130_fd_sc_hd__inv_2 _074_ (.A(net18),
    .Y(_027_));
 sky130_fd_sc_hd__inv_2 _075_ (.A(net18),
    .Y(_028_));
 sky130_fd_sc_hd__inv_2 _076_ (.A(net18),
    .Y(_029_));
 sky130_fd_sc_hd__inv_2 _077_ (.A(net18),
    .Y(_030_));
 sky130_fd_sc_hd__inv_2 _078_ (.A(net18),
    .Y(_031_));
 sky130_fd_sc_hd__dfrtp_1 _079_ (.CLK(clk),
    .D(\sine_out_temp[6] ),
    .RESET_B(_008_),
    .Q(net14));
 sky130_fd_sc_hd__dfrtp_1 _080_ (.CLK(clk),
    .D(\sine_out_temp[7] ),
    .RESET_B(_009_),
    .Q(net15));
 sky130_fd_sc_hd__dfrtp_1 _081_ (.CLK(clk),
    .D(\sine_out_temp[8] ),
    .RESET_B(_010_),
    .Q(net16));
 sky130_fd_sc_hd__dfrtp_1 _082_ (.CLK(clk),
    .D(\sine_out_temp[9] ),
    .RESET_B(_011_),
    .Q(net17));
 sky130_fd_sc_hd__dfrtp_1 _083_ (.CLK(clk),
    .D(\sine_out_temp[10] ),
    .RESET_B(_012_),
    .Q(net3));
 sky130_fd_sc_hd__dfrtp_1 _084_ (.CLK(clk),
    .D(\sine_out_temp[11] ),
    .RESET_B(_013_),
    .Q(net4));
 sky130_fd_sc_hd__dfrtp_1 _085_ (.CLK(clk),
    .D(\sine_out_temp[12] ),
    .RESET_B(_014_),
    .Q(net5));
 sky130_fd_sc_hd__dfrtp_1 _086_ (.CLK(clk),
    .D(\sine_out_temp[13] ),
    .RESET_B(_015_),
    .Q(net6));
 sky130_fd_sc_hd__dfrtp_1 _087_ (.CLK(clk),
    .D(\sine_out_temp[14] ),
    .RESET_B(_016_),
    .Q(net7));
 sky130_fd_sc_hd__dfrtp_1 _088_ (.CLK(clk),
    .D(\sine_out_temp[15] ),
    .RESET_B(_017_),
    .Q(net8));
 sky130_fd_sc_hd__dfrtp_4 _089_ (.CLK(clk),
    .D(_000_),
    .RESET_B(_018_),
    .Q(\tcout[0] ));
 sky130_fd_sc_hd__dfrtp_4 _090_ (.CLK(clk),
    .D(_001_),
    .RESET_B(_019_),
    .Q(\tcout[1] ));
 sky130_fd_sc_hd__dfrtp_1 _091_ (.CLK(clk),
    .D(_002_),
    .RESET_B(_020_),
    .Q(\tcout[2] ));
 sky130_fd_sc_hd__dfrtp_1 _092_ (.CLK(clk),
    .D(_003_),
    .RESET_B(_021_),
    .Q(\tcout[3] ));
 sky130_fd_sc_hd__dfrtp_1 _093_ (.CLK(clk),
    .D(_004_),
    .RESET_B(_022_),
    .Q(\tcout[4] ));
 sky130_fd_sc_hd__dfrtp_2 _094_ (.CLK(clk),
    .D(_005_),
    .RESET_B(_023_),
    .Q(\tcout[5] ));
 sky130_fd_sc_hd__dfrtp_1 _095_ (.CLK(clk),
    .D(_006_),
    .RESET_B(_024_),
    .Q(\tcout[6] ));
 sky130_fd_sc_hd__dfrtp_1 _096_ (.CLK(clk),
    .D(_007_),
    .RESET_B(_025_),
    .Q(\tcout[7] ));
 sky130_fd_sc_hd__dfrtp_1 _097_ (.CLK(clk),
    .D(\sine_out_temp[0] ),
    .RESET_B(_026_),
    .Q(net2));
 sky130_fd_sc_hd__dfrtp_1 _098_ (.CLK(clk),
    .D(\sine_out_temp[1] ),
    .RESET_B(_027_),
    .Q(net9));
 sky130_fd_sc_hd__dfrtp_1 _099_ (.CLK(clk),
    .D(\sine_out_temp[2] ),
    .RESET_B(_028_),
    .Q(net10));
 sky130_fd_sc_hd__dfrtp_1 _100_ (.CLK(clk),
    .D(\sine_out_temp[3] ),
    .RESET_B(_029_),
    .Q(net11));
 sky130_fd_sc_hd__dfrtp_1 _101_ (.CLK(clk),
    .D(\sine_out_temp[4] ),
    .RESET_B(_030_),
    .Q(net12));
 sky130_fd_sc_hd__dfrtp_1 _102_ (.CLK(clk),
    .D(\sine_out_temp[5] ),
    .RESET_B(_031_),
    .Q(net13));
 ram256x16 mem_i (.csb0(csb0),
    .csb1(net21),
    .clk0(clk),
    .clk1(clk),
    .addr0({addr0[7],
    addr0[6],
    addr0[5],
    addr0[4],
    addr0[3],
    addr0[2],
    addr0[1],
    addr0[0]}),
    .addr1({\tcout[7] ,
    \tcout[6] ,
    \tcout[5] ,
    \tcout[4] ,
    \tcout[3] ,
    \tcout[2] ,
    \tcout[1] ,
    \tcout[0] }),
    .din0({din0[15],
    din0[14],
    din0[13],
    din0[12],
    din0[11],
    din0[10],
    din0[9],
    din0[8],
    din0[7],
    din0[6],
    din0[5],
    din0[4],
    din0[3],
    din0[2],
    din0[1],
    din0[0]}),
    .dout1({\sine_out_temp[15] ,
    \sine_out_temp[14] ,
    \sine_out_temp[13] ,
    \sine_out_temp[12] ,
    \sine_out_temp[11] ,
    \sine_out_temp[10] ,
    \sine_out_temp[9] ,
    \sine_out_temp[8] ,
    \sine_out_temp[7] ,
    \sine_out_temp[6] ,
    \sine_out_temp[5] ,
    \sine_out_temp[4] ,
    \sine_out_temp[3] ,
    \sine_out_temp[2] ,
    \sine_out_temp[1] ,
    \sine_out_temp[0] }));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_117_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_118_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_119_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_120_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_121_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_122_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_123_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_124_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_125_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_126_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_127_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_2_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_2_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_2_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_2_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_2_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_2_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_2_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_2_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_2_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_2_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_2_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_2_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_2_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_2_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_2_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_2_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_2_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_2_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_2_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_2_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_2_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_2_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_2_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_2_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_2_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_2_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_2_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_2_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_2_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_2_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_2_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_2_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_2_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_2_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_2_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_2_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_2_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_2_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_2_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_2_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_2_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_2_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_2_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_2_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_2_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_2_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_2_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_2_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_2_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_2_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_2_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_2_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_2_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_2_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_2_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_2_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_2_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_2_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_2_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_2_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_2_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_2_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_2_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_2_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_2_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_2_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_2_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_2_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_2_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_2_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_2_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_2_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_2_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_2_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_2_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_2_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_2_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_2_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_2_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_2_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_2_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_2_Right_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_2_Right_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_2_Right_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_2_Right_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_2_Right_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_2_Right_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_2_Right_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_2_Right_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_2_Right_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_2_Right_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_2_Right_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_2_Right_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_2_Right_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_2_Right_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_2_Right_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_2_Right_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_2_Right_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_2_Right_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_2_Right_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_2_Right_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_2_Right_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_2_Right_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_2_Right_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_2_Right_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_2_Right_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_2_Right_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_1_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_1_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_1_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_1_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_1_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_1_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_1_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_1_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_1_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_1_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_1_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_1_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_1_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_1_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_1_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_1_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_1_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_1_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_1_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_1_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_1_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_1_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_1_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_1_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_1_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_1_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_1_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_1_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_1_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_1_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_1_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_1_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_1_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_1_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_1_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_1_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_1_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_1_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_1_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_1_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_1_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_1_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_1_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_1_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_1_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_1_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_1_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_1_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_1_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_1_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_1_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_1_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_1_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_1_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_1_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_1_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_1_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_1_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_1_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_1_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_1_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_1_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_1_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_1_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_1_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_1_Left_203 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_1_Left_204 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_1_Left_205 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_1_Left_206 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_1_Left_207 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_1_Left_208 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_1_Left_209 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_1_Left_210 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_1_Left_211 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_1_Left_212 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_1_Left_213 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_1_Left_214 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_1_Left_215 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_1_Left_216 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_1_Left_217 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_1_Left_218 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_1_Left_219 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_1_Left_220 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_1_Left_221 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_1_Left_222 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_1_Left_223 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_1_Left_224 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_1_Left_225 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_1_Left_226 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_1_Left_227 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_1_Left_228 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_1_Left_229 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_1_Left_230 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_1_Left_231 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_1_Left_232 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_1_Left_233 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_1_Left_234 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_1_Left_235 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_1_Left_236 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_1_Left_237 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_1_Left_238 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_1_Left_239 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_1_Left_240 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_1_Left_241 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_1_Left_242 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_1_Left_243 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_117_Left_244 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_118_Left_245 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_119_Left_246 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_120_Left_247 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_121_Left_248 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_122_Left_249 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_123_Left_250 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_124_Left_251 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_125_Left_252 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_126_Left_253 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_127_Left_254 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_1_Left_255 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_2_Left_256 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_2_Left_257 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_2_Left_258 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_2_Left_259 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_2_Left_260 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_2_Left_261 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_2_Left_262 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_2_Left_263 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_2_Left_264 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_2_Left_265 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_2_Left_266 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_2_Left_267 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_2_Left_268 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_2_Left_269 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_2_Left_270 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_2_Left_271 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_2_Left_272 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_2_Left_273 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_2_Left_274 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_2_Left_275 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_2_Left_276 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_2_Left_277 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_2_Left_278 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_2_Left_279 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_2_Left_280 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_2_Left_281 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_2_Left_282 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_2_Left_283 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_2_Left_284 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_2_Left_285 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_2_Left_286 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_2_Left_287 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_2_Left_288 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_2_Left_289 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_2_Left_290 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_2_Left_291 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_2_Left_292 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_2_Left_293 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_2_Left_294 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_2_Left_295 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_2_Left_296 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_2_Left_297 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_2_Left_298 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_2_Left_299 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_2_Left_300 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_2_Left_301 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_2_Left_302 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_2_Left_303 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_2_Left_304 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_2_Left_305 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_2_Left_306 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_2_Left_307 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_2_Left_308 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_2_Left_309 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_2_Left_310 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_2_Left_311 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_2_Left_312 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_2_Left_313 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_2_Left_314 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_2_Left_315 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_2_Left_316 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_2_Left_317 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_2_Left_318 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_2_Left_319 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_2_Left_320 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_2_Left_321 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_2_Left_322 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_2_Left_323 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_2_Left_324 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_2_Left_325 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_2_Left_326 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_2_Left_327 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_2_Left_328 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_2_Left_329 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_2_Left_330 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_2_Left_331 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_2_Left_332 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_2_Left_333 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_2_Left_334 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_2_Left_335 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_2_Left_336 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_2_Left_337 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_2_Left_338 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_2_Left_339 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_2_Left_340 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_2_Left_341 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_2_Left_342 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_2_Left_343 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_2_Left_344 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_2_Left_345 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_2_Left_346 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_2_Left_347 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_2_Left_348 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_2_Left_349 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_2_Left_350 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_2_Left_351 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_2_Left_352 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_2_Left_353 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_2_Left_354 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_2_Left_355 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_2_Left_356 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_2_Left_357 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_2_Left_358 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_2_Left_359 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_2_Left_360 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_2_Left_361 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_2_Left_362 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_1_Right_363 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_1_Right_364 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_1_Right_365 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_1_Right_366 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_1_Right_367 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_1_Right_368 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_1_Right_369 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_1_Right_370 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_1_Right_371 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_1_Right_372 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_1_Right_373 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_1_Right_374 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_1_Right_375 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_1_Right_376 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_1_Right_377 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_1_Right_378 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_1_Right_379 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_1_Right_380 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_1_Right_381 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_1_Right_382 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_1_Right_383 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_1_Right_384 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_1_Right_385 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_1_Right_386 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_1_Right_387 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_1_Right_388 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_1_Right_389 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_1_Right_390 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_1_Right_391 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_1_Right_392 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_1_Right_393 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_1_Right_394 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_1_Right_395 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_1_Right_396 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_1_Right_397 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_1_Right_398 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_1_Right_399 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_1_Right_400 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_1_Right_401 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_1_Right_402 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_1_Right_403 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_1_Right_404 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_1_Right_405 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_1_Right_406 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_1_Right_407 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_1_Right_408 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_1_Right_409 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_1_Right_410 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_1_Right_411 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_1_Right_412 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_1_Right_413 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_1_Right_414 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_1_Right_415 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_1_Right_416 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_1_Right_417 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_1_Right_418 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_1_Right_419 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_1_Right_420 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_1_Right_421 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_1_Right_422 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_1_Right_423 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_1_Right_424 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_1_Right_425 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_1_Right_426 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_1_Right_427 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_1_Right_428 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_1_Right_429 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_1_Right_430 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_1_Right_431 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_1_Right_432 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_1_Right_433 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_1_Right_434 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_1_Right_435 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_1_Right_436 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_1_Right_437 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_1_Right_438 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_1_Right_439 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_1_Right_440 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_1_Right_441 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_1_Right_442 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_1_Right_443 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_1_Right_444 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_1_Right_445 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_1_Right_446 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_1_Right_447 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_1_Right_448 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_1_Right_449 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_1_Right_450 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_1_Right_451 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_1_Right_452 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_1_Right_453 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_1_Right_454 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_1_Right_455 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_1_Right_456 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_1_Right_457 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_1_Right_458 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_1_Right_459 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_1_Right_460 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_1_Right_461 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_1_Right_462 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_1_Right_463 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_1_Right_464 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_1_Right_465 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_1_Right_466 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_1_Right_467 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_1_Right_468 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_1_Right_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_1_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_1_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_1_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_1_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_1_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_2_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_2_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_2_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_2_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_2_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_2_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_2_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_2_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_2_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_2_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_2_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_2_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_2_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_2_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_2_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_2_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_2_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_2_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_2_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_2_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_2_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_2_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_2_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_2_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_2_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_2_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_2_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_2_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_2_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_2_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_2_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_2_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_2_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_2_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_2_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_2_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_2_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_2_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_2_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_2_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_2_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_2_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_2_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_2_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_2_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_2_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_2_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_2_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_2_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_2_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_2_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_2_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_2_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_2_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_2_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_2_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2_1208 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(rst),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 output2 (.A(net2),
    .X(sine_out[0]));
 sky130_fd_sc_hd__clkbuf_1 output3 (.A(net3),
    .X(sine_out[10]));
 sky130_fd_sc_hd__clkbuf_1 output4 (.A(net4),
    .X(sine_out[11]));
 sky130_fd_sc_hd__clkbuf_1 output5 (.A(net5),
    .X(sine_out[12]));
 sky130_fd_sc_hd__clkbuf_1 output6 (.A(net6),
    .X(sine_out[13]));
 sky130_fd_sc_hd__clkbuf_1 output7 (.A(net7),
    .X(sine_out[14]));
 sky130_fd_sc_hd__clkbuf_1 output8 (.A(net8),
    .X(sine_out[15]));
 sky130_fd_sc_hd__clkbuf_1 output9 (.A(net9),
    .X(sine_out[1]));
 sky130_fd_sc_hd__clkbuf_1 output10 (.A(net10),
    .X(sine_out[2]));
 sky130_fd_sc_hd__clkbuf_1 output11 (.A(net11),
    .X(sine_out[3]));
 sky130_fd_sc_hd__clkbuf_1 output12 (.A(net12),
    .X(sine_out[4]));
 sky130_fd_sc_hd__clkbuf_1 output13 (.A(net13),
    .X(sine_out[5]));
 sky130_fd_sc_hd__clkbuf_1 output14 (.A(net14),
    .X(sine_out[6]));
 sky130_fd_sc_hd__clkbuf_1 output15 (.A(net15),
    .X(sine_out[7]));
 sky130_fd_sc_hd__clkbuf_1 output16 (.A(net16),
    .X(sine_out[8]));
 sky130_fd_sc_hd__clkbuf_1 output17 (.A(net17),
    .X(sine_out[9]));
 sky130_fd_sc_hd__buf_4 fanout18 (.A(net20),
    .X(net18));
 sky130_fd_sc_hd__buf_2 fanout19 (.A(net20),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_8 fanout20 (.A(net1),
    .X(net20));
 sky130_fd_sc_hd__conb_1 mem_i_21 (.LO(net21));
endmodule
