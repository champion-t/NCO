sine_table[0] = {
16'h0000,
16'h0218,
16'h0430,
16'h0648,
16'h085f,
16'h0a76,
16'h0c8c,
16'h0ea1,
16'h10b5,
16'h12c8,
16'h14da,
16'h16ea,
16'h18f9,
16'h1b05,
16'h1d11,
16'h1f1a,
16'h2121,
16'h2325,
16'h2528,
16'h2728,
16'h2925,
16'h2b1f,
16'h2d16,
16'h2f0a,
16'h30fb,
16'h32e9,
16'h34d3,
16'h36ba,
16'h389c,
16'h3a7b,
16'h3c56,
16'h3e2d,
16'h3fff,
16'h41ce,
16'h4397,
16'h455c,
16'h471c,
16'h48d8,
16'h4a8e,
16'h4c3f,
16'h4deb,
16'h4f92,
16'h5133,
16'h52cf,
16'h5465,
16'h55f5,
16'h577f,
16'h5904,
16'h5a82,
16'h5bfa,
16'h5d6b,
16'h5ed7,
16'h603c,
16'h619a,
16'h62f1,
16'h6442,
16'h658c,
16'h66cf,
16'h680b,
16'h693f,
16'h6a6d,
16'h6b93,
16'h6cb2,
16'h6dc9,
16'h6ed9,
16'h6fe1,
16'h70e2,
16'h71db,
16'h72cc,
16'h73b5,
16'h7496,
16'h7570,
16'h7641,
16'h770a,
16'h77cb,
16'h7884,
16'h7934,
16'h79dc,
16'h7a7c,
16'h7b13,
16'h7ba2,
16'h7c29,
16'h7ca7,
16'h7d1c,
16'h7d89,
16'h7dee,
16'h7e49,
16'h7e9c,
16'h7ee7,
16'h7f28,
16'h7f61,
16'h7f91,
16'h7fb9,
16'h7fd8,
16'h7fed,
16'h7ffb,
16'h7fff,
16'h7ffb,
16'h7fed,
16'h7fd8,
16'h7fb9,
16'h7f91,
16'h7f61,
16'h7f28,
16'h7ee7,
16'h7e9c,
16'h7e49,
16'h7dee,
16'h7d89,
16'h7d1c,
16'h7ca7,
16'h7c29,
16'h7ba2,
16'h7b13,
16'h7a7c,
16'h79dc,
16'h7934,
16'h7884,
16'h77cb,
16'h770a,
16'h7641,
16'h7570,
16'h7496,
16'h73b5,
16'h72cc,
16'h71db,
16'h70e2,
16'h6fe1,
16'h6ed9,
16'h6dc9,
16'h6cb2,
16'h6b93,
16'h6a6d,
16'h693f,
16'h680b,
16'h66cf,
16'h658c,
16'h6442,
16'h62f1,
16'h619a,
16'h603c,
16'h5ed7,
16'h5d6b,
16'h5bfa,
16'h5a82,
16'h5904,
16'h577f,
16'h55f5,
16'h5465,
16'h52cf,
16'h5133,
16'h4f92,
16'h4deb,
16'h4c3f,
16'h4a8e,
16'h48d8,
16'h471c,
16'h455c,
16'h4397,
16'h41ce,
16'h4000,
16'h3e2d,
16'h3c56,
16'h3a7b,
16'h389c,
16'h36ba,
16'h34d3,
16'h32e9,
16'h30fb,
16'h2f0a,
16'h2d16,
16'h2b1f,
16'h2925,
16'h2728,
16'h2528,
16'h2325,
16'h2121,
16'h1f1a,
16'h1d11,
16'h1b05,
16'h18f9,
16'h16ea,
16'h14da,
16'h12c8,
16'h10b5,
16'h0ea1,
16'h0c8c,
16'h0a76,
16'h085f,
16'h0648,
16'h0430,
16'h0218,
16'h0000,
16'hfde8,
16'hfbd0,
16'hf9b8,
16'hf7a1,
16'hf58a,
16'hf374,
16'hf15f,
16'hef4b,
16'hed38,
16'heb26,
16'he916,
16'he707,
16'he4fb,
16'he2ef,
16'he0e6,
16'hdedf,
16'hdcdb,
16'hdad8,
16'hd8d8,
16'hd6db,
16'hd4e1,
16'hd2ea,
16'hd0f6,
16'hcf05,
16'hcd17,
16'hcb2d,
16'hc946,
16'hc764,
16'hc585,
16'hc3aa,
16'hc1d3,
16'hc001,
16'hbe32,
16'hbc69,
16'hbaa4,
16'hb8e4,
16'hb728,
16'hb572,
16'hb3c1,
16'hb215,
16'hb06e,
16'haecd,
16'had31,
16'hab9b,
16'haa0b,
16'ha881,
16'ha6fc,
16'ha57e,
16'ha406,
16'ha295,
16'ha129,
16'h9fc4,
16'h9e66,
16'h9d0f,
16'h9bbe,
16'h9a74,
16'h9931,
16'h97f5,
16'h96c1,
16'h9593,
16'h946d,
16'h934e,
16'h9237
};