module counter (clk,
    rst,
    sine_out);
 input clk;
 input rst;
 output [15:0] sine_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire _369_;
 wire _370_;
 wire _371_;
 wire _372_;
 wire _373_;
 wire _374_;
 wire _375_;
 wire _376_;
 wire _377_;
 wire _378_;
 wire _379_;
 wire _380_;
 wire _381_;
 wire _382_;
 wire _383_;
 wire _384_;
 wire _385_;
 wire _386_;
 wire \tcout[0] ;
 wire \tcout[1] ;
 wire \tcout[2] ;
 wire \tcout[3] ;
 wire \tcout[4] ;
 wire \tcout[5] ;
 wire \tcout[6] ;
 wire \tcout[7] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;

 sky130_fd_sc_hd__inv_2 _387_ (.A(net79),
    .Y(_000_));
 sky130_fd_sc_hd__inv_2 _388_ (.A(net39),
    .Y(_328_));
 sky130_fd_sc_hd__inv_2 _389_ (.A(net43),
    .Y(_333_));
 sky130_fd_sc_hd__inv_2 _390_ (.A(net45),
    .Y(_334_));
 sky130_fd_sc_hd__inv_2 _391_ (.A(net56),
    .Y(_335_));
 sky130_fd_sc_hd__inv_2 _392_ (.A(net62),
    .Y(_336_));
 sky130_fd_sc_hd__inv_2 _393_ (.A(net35),
    .Y(_337_));
 sky130_fd_sc_hd__inv_2 _394_ (.A(net1),
    .Y(_008_));
 sky130_fd_sc_hd__nand2b_4 _395_ (.A_N(net73),
    .B(net56),
    .Y(_338_));
 sky130_fd_sc_hd__and2b_2 _396_ (.A_N(net63),
    .B(net53),
    .X(_339_));
 sky130_fd_sc_hd__nor2_2 _397_ (.A(net64),
    .B(net71),
    .Y(_340_));
 sky130_fd_sc_hd__or2_2 _398_ (.A(net65),
    .B(net73),
    .X(_341_));
 sky130_fd_sc_hd__nor3b_2 _399_ (.A(net65),
    .B(net73),
    .C_N(net56),
    .Y(_342_));
 sky130_fd_sc_hd__nand2_1 _400_ (.A(net54),
    .B(_340_),
    .Y(_343_));
 sky130_fd_sc_hd__and2b_1 _401_ (.A_N(net76),
    .B(net62),
    .X(_344_));
 sky130_fd_sc_hd__and2b_2 _402_ (.A_N(net65),
    .B(net78),
    .X(_345_));
 sky130_fd_sc_hd__nand2b_2 _403_ (.A_N(net61),
    .B(net75),
    .Y(_346_));
 sky130_fd_sc_hd__nand2_2 _404_ (.A(net78),
    .B(net66),
    .Y(_347_));
 sky130_fd_sc_hd__nor2_1 _405_ (.A(net76),
    .B(net63),
    .Y(_348_));
 sky130_fd_sc_hd__or2_2 _406_ (.A(net79),
    .B(net68),
    .X(_349_));
 sky130_fd_sc_hd__xnor2_4 _407_ (.A(net75),
    .B(net61),
    .Y(_350_));
 sky130_fd_sc_hd__nand2_1 _408_ (.A(net56),
    .B(_350_),
    .Y(_351_));
 sky130_fd_sc_hd__and2_1 _409_ (.A(net77),
    .B(net74),
    .X(_352_));
 sky130_fd_sc_hd__nand2_2 _410_ (.A(net75),
    .B(net70),
    .Y(_353_));
 sky130_fd_sc_hd__and3b_2 _411_ (.A_N(net65),
    .B(net74),
    .C(net78),
    .X(_354_));
 sky130_fd_sc_hd__a211o_1 _412_ (.A1(net59),
    .A2(_350_),
    .B1(_342_),
    .C1(net48),
    .X(_355_));
 sky130_fd_sc_hd__or2_2 _413_ (.A(net51),
    .B(net70),
    .X(_356_));
 sky130_fd_sc_hd__nand2_1 _414_ (.A(net27),
    .B(net67),
    .Y(_357_));
 sky130_fd_sc_hd__a21oi_1 _415_ (.A1(net74),
    .A2(_347_),
    .B1(net58),
    .Y(_358_));
 sky130_fd_sc_hd__nand2_2 _416_ (.A(net63),
    .B(net71),
    .Y(_359_));
 sky130_fd_sc_hd__and2b_1 _417_ (.A_N(net73),
    .B(net65),
    .X(_360_));
 sky130_fd_sc_hd__nand2b_2 _418_ (.A_N(net70),
    .B(net61),
    .Y(_361_));
 sky130_fd_sc_hd__nand2_1 _419_ (.A(net27),
    .B(_360_),
    .Y(_362_));
 sky130_fd_sc_hd__nand2_1 _420_ (.A(_346_),
    .B(_362_),
    .Y(_363_));
 sky130_fd_sc_hd__a2bb2o_1 _421_ (.A1_N(_355_),
    .A2_N(_358_),
    .B1(_363_),
    .B2(net49),
    .X(_364_));
 sky130_fd_sc_hd__nand2_1 _422_ (.A(net64),
    .B(net24),
    .Y(_365_));
 sky130_fd_sc_hd__and2b_1 _423_ (.A_N(net52),
    .B(net71),
    .X(_366_));
 sky130_fd_sc_hd__nand2b_1 _424_ (.A_N(net56),
    .B(net73),
    .Y(_367_));
 sky130_fd_sc_hd__o21bai_2 _425_ (.A1(net64),
    .A2(net71),
    .B1_N(net53),
    .Y(_368_));
 sky130_fd_sc_hd__a21o_1 _426_ (.A1(net67),
    .A2(net24),
    .B1(_368_),
    .X(_369_));
 sky130_fd_sc_hd__nand2_1 _427_ (.A(net76),
    .B(net54),
    .Y(_370_));
 sky130_fd_sc_hd__nand2_1 _428_ (.A(net58),
    .B(net24),
    .Y(_371_));
 sky130_fd_sc_hd__nor2_4 _429_ (.A(net32),
    .B(net49),
    .Y(_372_));
 sky130_fd_sc_hd__nand2b_1 _430_ (.A_N(net45),
    .B(net41),
    .Y(_373_));
 sky130_fd_sc_hd__or2_2 _431_ (.A(net77),
    .B(net74),
    .X(_374_));
 sky130_fd_sc_hd__xnor2_4 _432_ (.A(net75),
    .B(net70),
    .Y(_375_));
 sky130_fd_sc_hd__inv_2 _433_ (.A(_375_),
    .Y(_001_));
 sky130_fd_sc_hd__nor2_4 _434_ (.A(net32),
    .B(net29),
    .Y(_376_));
 sky130_fd_sc_hd__nand2_2 _435_ (.A(net41),
    .B(net45),
    .Y(_377_));
 sky130_fd_sc_hd__and2b_1 _436_ (.A_N(net78),
    .B(net73),
    .X(_378_));
 sky130_fd_sc_hd__nand2b_2 _437_ (.A_N(net78),
    .B(net73),
    .Y(_379_));
 sky130_fd_sc_hd__and2b_1 _438_ (.A_N(net63),
    .B(net71),
    .X(_380_));
 sky130_fd_sc_hd__nand2b_1 _439_ (.A_N(net67),
    .B(net74),
    .Y(_381_));
 sky130_fd_sc_hd__and2b_1 _440_ (.A_N(net72),
    .B(net75),
    .X(_382_));
 sky130_fd_sc_hd__nand2b_4 _441_ (.A_N(net74),
    .B(net77),
    .Y(_383_));
 sky130_fd_sc_hd__nand2_1 _442_ (.A(_339_),
    .B(_375_),
    .Y(_384_));
 sky130_fd_sc_hd__o311a_1 _443_ (.A1(net55),
    .A2(_344_),
    .A3(_354_),
    .B1(_384_),
    .C1(net48),
    .X(_385_));
 sky130_fd_sc_hd__a31o_1 _444_ (.A1(net31),
    .A2(_369_),
    .A3(_371_),
    .B1(_385_),
    .X(_386_));
 sky130_fd_sc_hd__mux2_1 _445_ (.A0(_364_),
    .A1(_386_),
    .S(net43),
    .X(_016_));
 sky130_fd_sc_hd__a21o_1 _446_ (.A1(_341_),
    .A2(_001_),
    .B1(net27),
    .X(_017_));
 sky130_fd_sc_hd__xnor2_4 _447_ (.A(net61),
    .B(net70),
    .Y(_018_));
 sky130_fd_sc_hd__nor2_1 _448_ (.A(_345_),
    .B(_018_),
    .Y(_019_));
 sky130_fd_sc_hd__o211ai_1 _449_ (.A1(net58),
    .A2(_019_),
    .B1(_017_),
    .C1(net49),
    .Y(_020_));
 sky130_fd_sc_hd__nor3_4 _450_ (.A(net76),
    .B(net64),
    .C(net71),
    .Y(_021_));
 sky130_fd_sc_hd__a21o_2 _451_ (.A1(net78),
    .A2(net66),
    .B1(net56),
    .X(_022_));
 sky130_fd_sc_hd__nand2_2 _452_ (.A(net51),
    .B(net70),
    .Y(_023_));
 sky130_fd_sc_hd__nand2_1 _453_ (.A(net56),
    .B(_378_),
    .Y(_024_));
 sky130_fd_sc_hd__and3_1 _454_ (.A(net52),
    .B(_353_),
    .C(_361_),
    .X(_025_));
 sky130_fd_sc_hd__nor2_1 _455_ (.A(net46),
    .B(_025_),
    .Y(_026_));
 sky130_fd_sc_hd__o21ai_1 _456_ (.A1(_021_),
    .A2(_022_),
    .B1(_026_),
    .Y(_027_));
 sky130_fd_sc_hd__nor2_1 _457_ (.A(net39),
    .B(net33),
    .Y(_028_));
 sky130_fd_sc_hd__nor2_2 _458_ (.A(net37),
    .B(net41),
    .Y(_029_));
 sky130_fd_sc_hd__or2_1 _459_ (.A(net37),
    .B(net42),
    .X(_030_));
 sky130_fd_sc_hd__a21boi_2 _460_ (.A1(net76),
    .A2(net69),
    .B1_N(net55),
    .Y(_031_));
 sky130_fd_sc_hd__a21bo_2 _461_ (.A1(net77),
    .A2(net67),
    .B1_N(net59),
    .X(_032_));
 sky130_fd_sc_hd__o311a_1 _462_ (.A1(_340_),
    .A2(_382_),
    .A3(_031_),
    .B1(_343_),
    .C1(net47),
    .X(_033_));
 sky130_fd_sc_hd__nand2_1 _463_ (.A(net58),
    .B(_019_),
    .Y(_034_));
 sky130_fd_sc_hd__and3b_1 _464_ (.A_N(net74),
    .B(net67),
    .C(net77),
    .X(_035_));
 sky130_fd_sc_hd__nand3b_1 _465_ (.A_N(net73),
    .B(net66),
    .C(net78),
    .Y(_036_));
 sky130_fd_sc_hd__nand2_1 _466_ (.A(net28),
    .B(_036_),
    .Y(_037_));
 sky130_fd_sc_hd__nor2_1 _467_ (.A(net50),
    .B(net57),
    .Y(_038_));
 sky130_fd_sc_hd__a31o_1 _468_ (.A1(net31),
    .A2(_034_),
    .A3(_037_),
    .B1(_033_),
    .X(_039_));
 sky130_fd_sc_hd__a32o_1 _469_ (.A1(_020_),
    .A2(_027_),
    .A3(_028_),
    .B1(_029_),
    .B2(_039_),
    .X(_040_));
 sky130_fd_sc_hd__o21bai_1 _470_ (.A1(net34),
    .A2(_016_),
    .B1_N(_040_),
    .Y(net2));
 sky130_fd_sc_hd__nor2_2 _471_ (.A(net51),
    .B(net62),
    .Y(_041_));
 sky130_fd_sc_hd__or2_1 _472_ (.A(net51),
    .B(net61),
    .X(_042_));
 sky130_fd_sc_hd__a221o_1 _473_ (.A1(_018_),
    .A2(_031_),
    .B1(_041_),
    .B2(net24),
    .C1(net30),
    .X(_043_));
 sky130_fd_sc_hd__and2_2 _474_ (.A(net59),
    .B(net67),
    .X(_044_));
 sky130_fd_sc_hd__nand2_2 _475_ (.A(net52),
    .B(net63),
    .Y(_045_));
 sky130_fd_sc_hd__nand2_1 _476_ (.A(net71),
    .B(_044_),
    .Y(_046_));
 sky130_fd_sc_hd__a32oi_1 _477_ (.A1(net76),
    .A2(_341_),
    .A3(_046_),
    .B1(_031_),
    .B2(net18),
    .Y(_047_));
 sky130_fd_sc_hd__o21ai_1 _478_ (.A1(net47),
    .A2(_047_),
    .B1(_043_),
    .Y(_048_));
 sky130_fd_sc_hd__nand2_1 _479_ (.A(net51),
    .B(_359_),
    .Y(_049_));
 sky130_fd_sc_hd__o21ai_1 _480_ (.A1(net75),
    .A2(net70),
    .B1(net61),
    .Y(_050_));
 sky130_fd_sc_hd__o21a_2 _481_ (.A1(net75),
    .A2(net70),
    .B1(net61),
    .X(_051_));
 sky130_fd_sc_hd__o21ai_2 _482_ (.A1(net76),
    .A2(net63),
    .B1(net53),
    .Y(_052_));
 sky130_fd_sc_hd__a2bb2o_1 _483_ (.A1_N(_051_),
    .A2_N(_052_),
    .B1(net26),
    .B2(_361_),
    .X(_053_));
 sky130_fd_sc_hd__nor2_1 _484_ (.A(_383_),
    .B(_045_),
    .Y(_054_));
 sky130_fd_sc_hd__and2b_2 _485_ (.A_N(net51),
    .B(net75),
    .X(_055_));
 sky130_fd_sc_hd__nand2_1 _486_ (.A(net66),
    .B(_353_),
    .Y(_056_));
 sky130_fd_sc_hd__a21boi_2 _487_ (.A1(net78),
    .A2(net74),
    .B1_N(net66),
    .Y(_057_));
 sky130_fd_sc_hd__a31o_1 _488_ (.A1(net75),
    .A2(net26),
    .A3(_018_),
    .B1(_054_),
    .X(_058_));
 sky130_fd_sc_hd__a221o_1 _489_ (.A1(_372_),
    .A2(_053_),
    .B1(_058_),
    .B2(_376_),
    .C1(net37),
    .X(_059_));
 sky130_fd_sc_hd__a21o_1 _490_ (.A1(net32),
    .A2(_048_),
    .B1(_059_),
    .X(_060_));
 sky130_fd_sc_hd__a21o_1 _491_ (.A1(net77),
    .A2(_018_),
    .B1(net27),
    .X(_061_));
 sky130_fd_sc_hd__nor2_1 _492_ (.A(net55),
    .B(_375_),
    .Y(_062_));
 sky130_fd_sc_hd__nand2_1 _493_ (.A(net26),
    .B(net18),
    .Y(_063_));
 sky130_fd_sc_hd__a31o_1 _494_ (.A1(_357_),
    .A2(_061_),
    .A3(_063_),
    .B1(net48),
    .X(_064_));
 sky130_fd_sc_hd__nand2_1 _495_ (.A(net65),
    .B(_379_),
    .Y(_065_));
 sky130_fd_sc_hd__o31a_1 _496_ (.A1(net57),
    .A2(_336_),
    .A3(_378_),
    .B1(net48),
    .X(_066_));
 sky130_fd_sc_hd__nand2_1 _497_ (.A(net55),
    .B(_374_),
    .Y(_067_));
 sky130_fd_sc_hd__o21ai_1 _498_ (.A1(_354_),
    .A2(_067_),
    .B1(_066_),
    .Y(_068_));
 sky130_fd_sc_hd__and3_1 _499_ (.A(net32),
    .B(_064_),
    .C(_068_),
    .X(_069_));
 sky130_fd_sc_hd__o32a_1 _500_ (.A1(net26),
    .A2(_345_),
    .A3(_382_),
    .B1(_356_),
    .B2(_350_),
    .X(_070_));
 sky130_fd_sc_hd__a21bo_1 _501_ (.A1(_338_),
    .A2(net23),
    .B1_N(_350_),
    .X(_071_));
 sky130_fd_sc_hd__a221o_1 _502_ (.A1(_376_),
    .A2(_070_),
    .B1(_071_),
    .B2(_372_),
    .C1(net34),
    .X(_072_));
 sky130_fd_sc_hd__o21a_1 _503_ (.A1(_069_),
    .A2(_072_),
    .B1(_337_),
    .X(_073_));
 sky130_fd_sc_hd__a221o_1 _504_ (.A1(net51),
    .A2(net70),
    .B1(_361_),
    .B2(_055_),
    .C1(_054_),
    .X(_074_));
 sky130_fd_sc_hd__a21o_1 _505_ (.A1(_347_),
    .A2(_349_),
    .B1(_049_),
    .X(_075_));
 sky130_fd_sc_hd__nor2_1 _506_ (.A(net48),
    .B(_055_),
    .Y(_076_));
 sky130_fd_sc_hd__a32o_1 _507_ (.A1(_362_),
    .A2(_075_),
    .A3(_076_),
    .B1(_074_),
    .B2(net44),
    .X(_077_));
 sky130_fd_sc_hd__a211o_2 _508_ (.A1(net76),
    .A2(net71),
    .B1(net63),
    .C1(net52),
    .X(_078_));
 sky130_fd_sc_hd__a21o_1 _509_ (.A1(_336_),
    .A2(_375_),
    .B1(_032_),
    .X(_079_));
 sky130_fd_sc_hd__a21o_1 _510_ (.A1(_078_),
    .A2(_079_),
    .B1(net22),
    .X(_080_));
 sky130_fd_sc_hd__a21oi_1 _511_ (.A1(net23),
    .A2(_042_),
    .B1(_350_),
    .Y(_081_));
 sky130_fd_sc_hd__o21ba_1 _512_ (.A1(_338_),
    .A2(_344_),
    .B1_N(_081_),
    .X(_082_));
 sky130_fd_sc_hd__o211a_1 _513_ (.A1(net21),
    .A2(_082_),
    .B1(_080_),
    .C1(net39),
    .X(_083_));
 sky130_fd_sc_hd__o21ai_1 _514_ (.A1(net41),
    .A2(_077_),
    .B1(_083_),
    .Y(_084_));
 sky130_fd_sc_hd__o211ai_1 _515_ (.A1(net56),
    .A2(_353_),
    .B1(_351_),
    .C1(net31),
    .Y(_085_));
 sky130_fd_sc_hd__or2_1 _516_ (.A(net77),
    .B(_368_),
    .X(_086_));
 sky130_fd_sc_hd__a31oi_1 _517_ (.A1(net49),
    .A2(_359_),
    .A3(_086_),
    .B1(net43),
    .Y(_087_));
 sky130_fd_sc_hd__nor2_1 _518_ (.A(net61),
    .B(_375_),
    .Y(_088_));
 sky130_fd_sc_hd__nand2_2 _519_ (.A(_336_),
    .B(_001_),
    .Y(_089_));
 sky130_fd_sc_hd__a21o_1 _520_ (.A1(_065_),
    .A2(_089_),
    .B1(net56),
    .X(_090_));
 sky130_fd_sc_hd__nor2_1 _521_ (.A(_347_),
    .B(net23),
    .Y(_091_));
 sky130_fd_sc_hd__a31o_1 _522_ (.A1(_347_),
    .A2(net23),
    .A3(_383_),
    .B1(_091_),
    .X(_092_));
 sky130_fd_sc_hd__a221o_1 _523_ (.A1(_085_),
    .A2(_087_),
    .B1(_092_),
    .B2(_372_),
    .C1(net39),
    .X(_093_));
 sky130_fd_sc_hd__a31o_1 _524_ (.A1(_376_),
    .A2(_024_),
    .A3(_090_),
    .B1(_093_),
    .X(_094_));
 sky130_fd_sc_hd__a32o_1 _525_ (.A1(net35),
    .A2(_084_),
    .A3(_094_),
    .B1(_060_),
    .B2(_073_),
    .X(net9));
 sky130_fd_sc_hd__o21ai_1 _526_ (.A1(net65),
    .A2(net73),
    .B1(net57),
    .Y(_095_));
 sky130_fd_sc_hd__a21oi_1 _527_ (.A1(net65),
    .A2(net18),
    .B1(_095_),
    .Y(_096_));
 sky130_fd_sc_hd__a211oi_1 _528_ (.A1(_341_),
    .A2(_062_),
    .B1(_096_),
    .C1(net22),
    .Y(_097_));
 sky130_fd_sc_hd__nor3b_1 _529_ (.A(net78),
    .B(net66),
    .C_N(net73),
    .Y(_098_));
 sky130_fd_sc_hd__nor2_1 _530_ (.A(_336_),
    .B(_382_),
    .Y(_099_));
 sky130_fd_sc_hd__or3_1 _531_ (.A(net57),
    .B(_035_),
    .C(_098_),
    .X(_100_));
 sky130_fd_sc_hd__nand2_1 _532_ (.A(_379_),
    .B(_044_),
    .Y(_101_));
 sky130_fd_sc_hd__a21oi_2 _533_ (.A1(_379_),
    .A2(_044_),
    .B1(net31),
    .Y(_102_));
 sky130_fd_sc_hd__a221oi_1 _534_ (.A1(_038_),
    .A2(_056_),
    .B1(_100_),
    .B2(_102_),
    .C1(\tcout[5] ),
    .Y(_103_));
 sky130_fd_sc_hd__o211a_1 _535_ (.A1(_018_),
    .A2(_022_),
    .B1(_024_),
    .C1(_376_),
    .X(_104_));
 sky130_fd_sc_hd__or4_1 _536_ (.A(net34),
    .B(_097_),
    .C(_103_),
    .D(_104_),
    .X(_105_));
 sky130_fd_sc_hd__nor2_1 _537_ (.A(_378_),
    .B(_022_),
    .Y(_106_));
 sky130_fd_sc_hd__a21oi_1 _538_ (.A1(_065_),
    .A2(_089_),
    .B1(net27),
    .Y(_107_));
 sky130_fd_sc_hd__o21a_1 _539_ (.A1(_106_),
    .A2(_107_),
    .B1(_372_),
    .X(_108_));
 sky130_fd_sc_hd__o211a_1 _540_ (.A1(net27),
    .A2(_057_),
    .B1(_076_),
    .C1(_362_),
    .X(_109_));
 sky130_fd_sc_hd__o311a_1 _541_ (.A1(_339_),
    .A2(_344_),
    .A3(_382_),
    .B1(_338_),
    .C1(net44),
    .X(_110_));
 sky130_fd_sc_hd__a31o_1 _542_ (.A1(net57),
    .A2(_374_),
    .A3(_381_),
    .B1(net21),
    .X(_111_));
 sky130_fd_sc_hd__o31ai_1 _543_ (.A1(net43),
    .A2(_109_),
    .A3(_110_),
    .B1(_111_),
    .Y(_112_));
 sky130_fd_sc_hd__o311a_1 _544_ (.A1(net39),
    .A2(_108_),
    .A3(_112_),
    .B1(net35),
    .C1(_105_),
    .X(_113_));
 sky130_fd_sc_hd__a21oi_1 _545_ (.A1(net27),
    .A2(_019_),
    .B1(_355_),
    .Y(_114_));
 sky130_fd_sc_hd__and3b_1 _546_ (.A_N(net53),
    .B(net63),
    .C(net72),
    .X(_115_));
 sky130_fd_sc_hd__nand3b_1 _547_ (.A_N(net52),
    .B(net64),
    .C(net71),
    .Y(_116_));
 sky130_fd_sc_hd__o311a_1 _548_ (.A1(_366_),
    .A2(_025_),
    .A3(_055_),
    .B1(_116_),
    .C1(net46),
    .X(_117_));
 sky130_fd_sc_hd__o21a_1 _549_ (.A1(_114_),
    .A2(_117_),
    .B1(net32),
    .X(_118_));
 sky130_fd_sc_hd__o221a_1 _550_ (.A1(net77),
    .A2(_359_),
    .B1(_383_),
    .B2(net67),
    .C1(net58),
    .X(_119_));
 sky130_fd_sc_hd__nor2_1 _551_ (.A(net58),
    .B(_345_),
    .Y(_120_));
 sky130_fd_sc_hd__a21o_1 _552_ (.A1(_374_),
    .A2(_120_),
    .B1(_119_),
    .X(_121_));
 sky130_fd_sc_hd__nand2_4 _553_ (.A(net62),
    .B(_375_),
    .Y(_122_));
 sky130_fd_sc_hd__nand2_1 _554_ (.A(net23),
    .B(_122_),
    .Y(_123_));
 sky130_fd_sc_hd__a32o_1 _555_ (.A1(_357_),
    .A2(_376_),
    .A3(_123_),
    .B1(_121_),
    .B2(_372_),
    .X(_124_));
 sky130_fd_sc_hd__or3_1 _556_ (.A(net34),
    .B(_118_),
    .C(_124_),
    .X(_125_));
 sky130_fd_sc_hd__a21o_1 _557_ (.A1(_336_),
    .A2(_375_),
    .B1(_051_),
    .X(_126_));
 sky130_fd_sc_hd__a31o_1 _558_ (.A1(_349_),
    .A2(_381_),
    .A3(_036_),
    .B1(net57),
    .X(_127_));
 sky130_fd_sc_hd__nor2_1 _559_ (.A(_349_),
    .B(net23),
    .Y(_128_));
 sky130_fd_sc_hd__a21o_1 _560_ (.A1(_126_),
    .A2(_127_),
    .B1(_128_),
    .X(_129_));
 sky130_fd_sc_hd__o221a_1 _561_ (.A1(net57),
    .A2(_019_),
    .B1(_032_),
    .B2(_088_),
    .C1(net48),
    .X(_130_));
 sky130_fd_sc_hd__or3_1 _562_ (.A(net39),
    .B(net32),
    .C(_130_),
    .X(_131_));
 sky130_fd_sc_hd__o22a_1 _563_ (.A1(_350_),
    .A2(_356_),
    .B1(_375_),
    .B2(_045_),
    .X(_132_));
 sky130_fd_sc_hd__nor2_1 _564_ (.A(net47),
    .B(_132_),
    .Y(_133_));
 sky130_fd_sc_hd__o21ai_2 _565_ (.A1(_366_),
    .A2(_041_),
    .B1(_350_),
    .Y(_134_));
 sky130_fd_sc_hd__a211o_1 _566_ (.A1(_102_),
    .A2(_134_),
    .B1(_133_),
    .C1(net20),
    .X(_135_));
 sky130_fd_sc_hd__a22o_1 _567_ (.A1(_372_),
    .A2(_129_),
    .B1(_131_),
    .B2(_135_),
    .X(_136_));
 sky130_fd_sc_hd__a31o_1 _568_ (.A1(_337_),
    .A2(_125_),
    .A3(_136_),
    .B1(_113_),
    .X(net10));
 sky130_fd_sc_hd__nor3b_1 _569_ (.A(net77),
    .B(\tcout[1] ),
    .C_N(net67),
    .Y(_137_));
 sky130_fd_sc_hd__nor3_1 _570_ (.A(net58),
    .B(_345_),
    .C(net19),
    .Y(_138_));
 sky130_fd_sc_hd__o21a_1 _571_ (.A1(_119_),
    .A2(_138_),
    .B1(net31),
    .X(_139_));
 sky130_fd_sc_hd__a21o_1 _572_ (.A1(net67),
    .A2(_001_),
    .B1(net58),
    .X(_140_));
 sky130_fd_sc_hd__or2_1 _573_ (.A(_380_),
    .B(_052_),
    .X(_141_));
 sky130_fd_sc_hd__o211a_1 _574_ (.A1(_035_),
    .A2(_141_),
    .B1(_140_),
    .C1(net49),
    .X(_142_));
 sky130_fd_sc_hd__o21a_1 _575_ (.A1(_139_),
    .A2(_142_),
    .B1(net33),
    .X(_143_));
 sky130_fd_sc_hd__nand2_1 _576_ (.A(_383_),
    .B(_120_),
    .Y(_144_));
 sky130_fd_sc_hd__a21oi_1 _577_ (.A1(_061_),
    .A2(_144_),
    .B1(net21),
    .Y(_145_));
 sky130_fd_sc_hd__a211o_1 _578_ (.A1(net69),
    .A2(net18),
    .B1(_354_),
    .C1(net58),
    .X(_146_));
 sky130_fd_sc_hd__nor2_1 _579_ (.A(_340_),
    .B(_052_),
    .Y(_147_));
 sky130_fd_sc_hd__or3_2 _580_ (.A(_340_),
    .B(_051_),
    .C(_052_),
    .X(_148_));
 sky130_fd_sc_hd__and3_1 _581_ (.A(_372_),
    .B(_146_),
    .C(_148_),
    .X(_149_));
 sky130_fd_sc_hd__or4_1 _582_ (.A(net34),
    .B(_143_),
    .C(_145_),
    .D(_149_),
    .X(_150_));
 sky130_fd_sc_hd__o21ai_1 _583_ (.A1(_035_),
    .A2(_141_),
    .B1(_362_),
    .Y(_151_));
 sky130_fd_sc_hd__o211a_1 _584_ (.A1(_352_),
    .A2(_032_),
    .B1(_369_),
    .C1(net31),
    .X(_152_));
 sky130_fd_sc_hd__a211o_1 _585_ (.A1(net49),
    .A2(_151_),
    .B1(_152_),
    .C1(net43),
    .X(_153_));
 sky130_fd_sc_hd__a221o_1 _586_ (.A1(_102_),
    .A2(_134_),
    .B1(_141_),
    .B2(_146_),
    .C1(net39),
    .X(_154_));
 sky130_fd_sc_hd__nand2_1 _587_ (.A(net20),
    .B(_154_),
    .Y(_155_));
 sky130_fd_sc_hd__a21oi_1 _588_ (.A1(_153_),
    .A2(_155_),
    .B1(net36),
    .Y(_156_));
 sky130_fd_sc_hd__a21oi_2 _589_ (.A1(net63),
    .A2(net72),
    .B1(net53),
    .Y(_157_));
 sky130_fd_sc_hd__nand2_1 _590_ (.A(_089_),
    .B(_157_),
    .Y(_158_));
 sky130_fd_sc_hd__a221o_1 _591_ (.A1(net46),
    .A2(_151_),
    .B1(_158_),
    .B2(_026_),
    .C1(net42),
    .X(_159_));
 sky130_fd_sc_hd__o311a_1 _592_ (.A1(net46),
    .A2(net71),
    .A3(_348_),
    .B1(_045_),
    .C1(net42),
    .X(_160_));
 sky130_fd_sc_hd__nand2_1 _593_ (.A(_134_),
    .B(_160_),
    .Y(_161_));
 sky130_fd_sc_hd__a21o_1 _594_ (.A1(_159_),
    .A2(_161_),
    .B1(net39),
    .X(_162_));
 sky130_fd_sc_hd__o21ai_1 _595_ (.A1(_035_),
    .A2(_052_),
    .B1(_140_),
    .Y(_163_));
 sky130_fd_sc_hd__a21oi_1 _596_ (.A1(_146_),
    .A2(_148_),
    .B1(net22),
    .Y(_164_));
 sky130_fd_sc_hd__and2_1 _597_ (.A(_339_),
    .B(_353_),
    .X(_165_));
 sky130_fd_sc_hd__nand2_1 _598_ (.A(_339_),
    .B(net18),
    .Y(_166_));
 sky130_fd_sc_hd__nand2_1 _599_ (.A(_349_),
    .B(_157_),
    .Y(_167_));
 sky130_fd_sc_hd__a31o_1 _600_ (.A1(_046_),
    .A2(_166_),
    .A3(_167_),
    .B1(net21),
    .X(_168_));
 sky130_fd_sc_hd__or3b_1 _601_ (.A(net34),
    .B(_164_),
    .C_N(_168_),
    .X(_169_));
 sky130_fd_sc_hd__a31o_1 _602_ (.A1(net33),
    .A2(_027_),
    .A3(_163_),
    .B1(_169_),
    .X(_170_));
 sky130_fd_sc_hd__a32o_1 _603_ (.A1(net36),
    .A2(_162_),
    .A3(_170_),
    .B1(_150_),
    .B2(_156_),
    .X(net11));
 sky130_fd_sc_hd__nor2_1 _604_ (.A(net45),
    .B(_115_),
    .Y(_171_));
 sky130_fd_sc_hd__and3_1 _605_ (.A(net29),
    .B(_078_),
    .C(_116_),
    .X(_172_));
 sky130_fd_sc_hd__a21o_1 _606_ (.A1(net63),
    .A2(_383_),
    .B1(_368_),
    .X(_173_));
 sky130_fd_sc_hd__a21oi_1 _607_ (.A1(_383_),
    .A2(_044_),
    .B1(net29),
    .Y(_174_));
 sky130_fd_sc_hd__a22oi_1 _608_ (.A1(_148_),
    .A2(_172_),
    .B1(_173_),
    .B2(_174_),
    .Y(_175_));
 sky130_fd_sc_hd__nor2_1 _609_ (.A(_380_),
    .B(_032_),
    .Y(_176_));
 sky130_fd_sc_hd__o2111a_1 _610_ (.A1(_380_),
    .A2(_032_),
    .B1(net42),
    .C1(_353_),
    .D1(_368_),
    .X(_177_));
 sky130_fd_sc_hd__and3_1 _611_ (.A(net44),
    .B(_353_),
    .C(_361_),
    .X(_178_));
 sky130_fd_sc_hd__o31ai_4 _612_ (.A1(net75),
    .A2(net61),
    .A3(net70),
    .B1(net51),
    .Y(_179_));
 sky130_fd_sc_hd__a2bb2o_1 _613_ (.A1_N(_376_),
    .A2_N(_177_),
    .B1(_178_),
    .B2(_179_),
    .X(_180_));
 sky130_fd_sc_hd__o211a_1 _614_ (.A1(net41),
    .A2(_175_),
    .B1(_180_),
    .C1(net37),
    .X(_181_));
 sky130_fd_sc_hd__o211a_1 _615_ (.A1(net62),
    .A2(net18),
    .B1(_050_),
    .C1(net26),
    .X(_182_));
 sky130_fd_sc_hd__a211o_1 _616_ (.A1(_122_),
    .A2(_147_),
    .B1(_182_),
    .C1(net22),
    .X(_183_));
 sky130_fd_sc_hd__o211ai_2 _617_ (.A1(net61),
    .A2(_375_),
    .B1(_359_),
    .C1(net51),
    .Y(_184_));
 sky130_fd_sc_hd__a31o_1 _618_ (.A1(net23),
    .A2(_042_),
    .A3(_184_),
    .B1(net21),
    .X(_185_));
 sky130_fd_sc_hd__and3_1 _619_ (.A(net34),
    .B(_183_),
    .C(_185_),
    .X(_186_));
 sky130_fd_sc_hd__nand4_1 _620_ (.A(_338_),
    .B(_032_),
    .C(_066_),
    .D(_078_),
    .Y(_187_));
 sky130_fd_sc_hd__a31o_1 _621_ (.A1(net51),
    .A2(_346_),
    .A3(_361_),
    .B1(net44),
    .X(_188_));
 sky130_fd_sc_hd__a21o_1 _622_ (.A1(_187_),
    .A2(_188_),
    .B1(net41),
    .X(_189_));
 sky130_fd_sc_hd__a21oi_1 _623_ (.A1(_186_),
    .A2(_189_),
    .B1(_181_),
    .Y(_190_));
 sky130_fd_sc_hd__a31o_1 _624_ (.A1(_346_),
    .A2(_361_),
    .A3(net23),
    .B1(net44),
    .X(_191_));
 sky130_fd_sc_hd__a21o_1 _625_ (.A1(_187_),
    .A2(_191_),
    .B1(net20),
    .X(_192_));
 sky130_fd_sc_hd__o211a_1 _626_ (.A1(_181_),
    .A2(_186_),
    .B1(_192_),
    .C1(net35),
    .X(_193_));
 sky130_fd_sc_hd__a21oi_1 _627_ (.A1(net25),
    .A2(_190_),
    .B1(_193_),
    .Y(net12));
 sky130_fd_sc_hd__o211ai_1 _628_ (.A1(_021_),
    .A2(_032_),
    .B1(_134_),
    .C1(net46),
    .Y(_194_));
 sky130_fd_sc_hd__nand2_1 _629_ (.A(_076_),
    .B(_184_),
    .Y(_195_));
 sky130_fd_sc_hd__a21oi_1 _630_ (.A1(_194_),
    .A2(_195_),
    .B1(net20),
    .Y(_196_));
 sky130_fd_sc_hd__and4_1 _631_ (.A(net28),
    .B(_349_),
    .C(_381_),
    .D(_036_),
    .X(_197_));
 sky130_fd_sc_hd__nand2_1 _632_ (.A(_028_),
    .B(_102_),
    .Y(_198_));
 sky130_fd_sc_hd__nor2_1 _633_ (.A(net37),
    .B(_373_),
    .Y(_199_));
 sky130_fd_sc_hd__or4b_1 _634_ (.A(_055_),
    .B(net19),
    .C(_176_),
    .D_N(_199_),
    .X(_200_));
 sky130_fd_sc_hd__o21ai_1 _635_ (.A1(_197_),
    .A2(_198_),
    .B1(_200_),
    .Y(_201_));
 sky130_fd_sc_hd__a32o_1 _636_ (.A1(net54),
    .A2(_089_),
    .A3(_122_),
    .B1(_120_),
    .B2(_374_),
    .X(_202_));
 sky130_fd_sc_hd__o211a_1 _637_ (.A1(_349_),
    .A2(net23),
    .B1(net46),
    .C1(_338_),
    .X(_203_));
 sky130_fd_sc_hd__a31o_1 _638_ (.A1(_370_),
    .A2(_122_),
    .A3(_203_),
    .B1(net41),
    .X(_204_));
 sky130_fd_sc_hd__a21o_1 _639_ (.A1(net30),
    .A2(_202_),
    .B1(_204_),
    .X(_205_));
 sky130_fd_sc_hd__and2_1 _640_ (.A(_343_),
    .B(_370_),
    .X(_206_));
 sky130_fd_sc_hd__nand2_1 _641_ (.A(net77),
    .B(_342_),
    .Y(_207_));
 sky130_fd_sc_hd__o2111a_1 _642_ (.A1(_339_),
    .A2(_379_),
    .B1(_207_),
    .C1(_357_),
    .D1(net29),
    .X(_208_));
 sky130_fd_sc_hd__a311o_1 _643_ (.A1(net46),
    .A2(_158_),
    .A3(_206_),
    .B1(_208_),
    .C1(net32),
    .X(_209_));
 sky130_fd_sc_hd__a31o_1 _644_ (.A1(net38),
    .A2(_205_),
    .A3(_209_),
    .B1(_201_),
    .X(_210_));
 sky130_fd_sc_hd__a311o_1 _645_ (.A1(net38),
    .A2(_205_),
    .A3(_209_),
    .B1(_196_),
    .C1(_201_),
    .X(_211_));
 sky130_fd_sc_hd__a31o_1 _646_ (.A1(_046_),
    .A2(_086_),
    .A3(_166_),
    .B1(net46),
    .X(_212_));
 sky130_fd_sc_hd__a21o_1 _647_ (.A1(_194_),
    .A2(_212_),
    .B1(net20),
    .X(_213_));
 sky130_fd_sc_hd__nand2_1 _648_ (.A(net35),
    .B(_213_),
    .Y(_214_));
 sky130_fd_sc_hd__o2bb2a_1 _649_ (.A1_N(net25),
    .A2_N(_211_),
    .B1(_214_),
    .B2(_210_),
    .X(net13));
 sky130_fd_sc_hd__a221o_1 _650_ (.A1(net24),
    .A2(_041_),
    .B1(_051_),
    .B2(net26),
    .C1(net45),
    .X(_215_));
 sky130_fd_sc_hd__a31oi_1 _651_ (.A1(net52),
    .A2(_346_),
    .A3(_122_),
    .B1(_215_),
    .Y(_216_));
 sky130_fd_sc_hd__nand2_1 _652_ (.A(net18),
    .B(_041_),
    .Y(_217_));
 sky130_fd_sc_hd__a41o_1 _653_ (.A1(net44),
    .A2(_365_),
    .A3(_207_),
    .A4(_217_),
    .B1(net41),
    .X(_218_));
 sky130_fd_sc_hd__nor2_1 _654_ (.A(_340_),
    .B(net18),
    .Y(_219_));
 sky130_fd_sc_hd__nor2_1 _655_ (.A(net52),
    .B(_021_),
    .Y(_220_));
 sky130_fd_sc_hd__o21ai_1 _656_ (.A1(_219_),
    .A2(_220_),
    .B1(_376_),
    .Y(_221_));
 sky130_fd_sc_hd__a21oi_1 _657_ (.A1(_089_),
    .A2(_122_),
    .B1(net27),
    .Y(_222_));
 sky130_fd_sc_hd__o211ai_1 _658_ (.A1(net28),
    .A2(_122_),
    .B1(_089_),
    .C1(_372_),
    .Y(_223_));
 sky130_fd_sc_hd__o211ai_1 _659_ (.A1(_216_),
    .A2(_218_),
    .B1(_221_),
    .C1(_223_),
    .Y(_224_));
 sky130_fd_sc_hd__o211a_1 _660_ (.A1(net67),
    .A2(_383_),
    .B1(_359_),
    .C1(net59),
    .X(_225_));
 sky130_fd_sc_hd__or3b_1 _661_ (.A(net22),
    .B(_225_),
    .C_N(_369_),
    .X(_226_));
 sky130_fd_sc_hd__a211o_1 _662_ (.A1(_383_),
    .A2(_044_),
    .B1(_358_),
    .C1(_377_),
    .X(_227_));
 sky130_fd_sc_hd__a21oi_1 _663_ (.A1(_226_),
    .A2(_227_),
    .B1(net39),
    .Y(_228_));
 sky130_fd_sc_hd__a21o_1 _664_ (.A1(_049_),
    .A2(_173_),
    .B1(net29),
    .X(_229_));
 sky130_fd_sc_hd__a21o_1 _665_ (.A1(_356_),
    .A2(_179_),
    .B1(net44),
    .X(_230_));
 sky130_fd_sc_hd__a21oi_1 _666_ (.A1(_229_),
    .A2(_230_),
    .B1(net20),
    .Y(_231_));
 sky130_fd_sc_hd__a211oi_1 _667_ (.A1(net37),
    .A2(_224_),
    .B1(_228_),
    .C1(_231_),
    .Y(_232_));
 sky130_fd_sc_hd__o31ai_1 _668_ (.A1(net45),
    .A2(_366_),
    .A3(_021_),
    .B1(_229_),
    .Y(_233_));
 sky130_fd_sc_hd__a221o_1 _669_ (.A1(net37),
    .A2(_224_),
    .B1(_233_),
    .B2(_029_),
    .C1(_228_),
    .X(_234_));
 sky130_fd_sc_hd__mux2_1 _670_ (.A0(_232_),
    .A1(_234_),
    .S(net35),
    .X(net14));
 sky130_fd_sc_hd__a31o_1 _671_ (.A1(net27),
    .A2(net65),
    .A3(_379_),
    .B1(net50),
    .X(_235_));
 sky130_fd_sc_hd__o32a_1 _672_ (.A1(_334_),
    .A2(_021_),
    .A3(_055_),
    .B1(_096_),
    .B2(_235_),
    .X(_236_));
 sky130_fd_sc_hd__o31ai_1 _673_ (.A1(net21),
    .A2(_051_),
    .A3(_220_),
    .B1(net37),
    .Y(_237_));
 sky130_fd_sc_hd__a21oi_1 _674_ (.A1(_336_),
    .A2(_383_),
    .B1(_022_),
    .Y(_238_));
 sky130_fd_sc_hd__a21o_1 _675_ (.A1(_379_),
    .A2(_031_),
    .B1(net22),
    .X(_239_));
 sky130_fd_sc_hd__o22ai_1 _676_ (.A1(net43),
    .A2(_236_),
    .B1(_238_),
    .B2(_239_),
    .Y(_240_));
 sky130_fd_sc_hd__a2111o_1 _677_ (.A1(net72),
    .A2(_344_),
    .B1(_345_),
    .C1(_382_),
    .D1(net26),
    .X(_241_));
 sky130_fd_sc_hd__a32o_1 _678_ (.A1(net29),
    .A2(_042_),
    .A3(_179_),
    .B1(_241_),
    .B2(_066_),
    .X(_242_));
 sky130_fd_sc_hd__and2_1 _679_ (.A(net32),
    .B(_242_),
    .X(_243_));
 sky130_fd_sc_hd__or3_1 _680_ (.A(net52),
    .B(net24),
    .C(_380_),
    .X(_244_));
 sky130_fd_sc_hd__o21a_1 _681_ (.A1(_051_),
    .A2(_052_),
    .B1(_376_),
    .X(_245_));
 sky130_fd_sc_hd__a221o_1 _682_ (.A1(_372_),
    .A2(_206_),
    .B1(_244_),
    .B2(_245_),
    .C1(net38),
    .X(_246_));
 sky130_fd_sc_hd__o22a_1 _683_ (.A1(_237_),
    .A2(_240_),
    .B1(_243_),
    .B2(_246_),
    .X(_247_));
 sky130_fd_sc_hd__nand2_1 _684_ (.A(_021_),
    .B(_038_),
    .Y(_248_));
 sky130_fd_sc_hd__and2_1 _685_ (.A(net35),
    .B(_248_),
    .X(_249_));
 sky130_fd_sc_hd__mux2_1 _686_ (.A0(_249_),
    .A1(net25),
    .S(_247_),
    .X(net15));
 sky130_fd_sc_hd__o21ai_1 _687_ (.A1(net49),
    .A2(_023_),
    .B1(_028_),
    .Y(_250_));
 sky130_fd_sc_hd__a31o_1 _688_ (.A1(net49),
    .A2(_144_),
    .A3(_166_),
    .B1(_250_),
    .X(_251_));
 sky130_fd_sc_hd__a22o_1 _689_ (.A1(net44),
    .A2(_062_),
    .B1(_079_),
    .B2(_171_),
    .X(_252_));
 sky130_fd_sc_hd__o21a_1 _690_ (.A1(net76),
    .A2(_368_),
    .B1(_370_),
    .X(_253_));
 sky130_fd_sc_hd__o21ai_1 _691_ (.A1(net21),
    .A2(_253_),
    .B1(net38),
    .Y(_254_));
 sky130_fd_sc_hd__or3_1 _692_ (.A(net26),
    .B(_350_),
    .C(net24),
    .X(_255_));
 sky130_fd_sc_hd__o211a_1 _693_ (.A1(net19),
    .A2(_244_),
    .B1(_255_),
    .C1(_372_),
    .X(_256_));
 sky130_fd_sc_hd__a211o_1 _694_ (.A1(net33),
    .A2(_252_),
    .B1(_254_),
    .C1(_256_),
    .X(_257_));
 sky130_fd_sc_hd__nand2_1 _695_ (.A(_251_),
    .B(_257_),
    .Y(_258_));
 sky130_fd_sc_hd__o21ai_1 _696_ (.A1(net58),
    .A2(_374_),
    .B1(_381_),
    .Y(_259_));
 sky130_fd_sc_hd__o221a_1 _697_ (.A1(_346_),
    .A2(net23),
    .B1(_259_),
    .B2(net24),
    .C1(net49),
    .X(_260_));
 sky130_fd_sc_hd__a21oi_1 _698_ (.A1(_086_),
    .A2(_206_),
    .B1(net46),
    .Y(_261_));
 sky130_fd_sc_hd__o21a_1 _699_ (.A1(_260_),
    .A2(_261_),
    .B1(_029_),
    .X(_262_));
 sky130_fd_sc_hd__o21a_1 _700_ (.A1(net78),
    .A2(_095_),
    .B1(_076_),
    .X(_263_));
 sky130_fd_sc_hd__o21ai_1 _701_ (.A1(_260_),
    .A2(_263_),
    .B1(_029_),
    .Y(_264_));
 sky130_fd_sc_hd__a31o_1 _702_ (.A1(_251_),
    .A2(_257_),
    .A3(_264_),
    .B1(net36),
    .X(_265_));
 sky130_fd_sc_hd__o31a_1 _703_ (.A1(net25),
    .A2(_258_),
    .A3(_262_),
    .B1(_265_),
    .X(net16));
 sky130_fd_sc_hd__a21o_1 _704_ (.A1(net79),
    .A2(net52),
    .B1(_197_),
    .X(_266_));
 sky130_fd_sc_hd__o211a_1 _705_ (.A1(_340_),
    .A2(net18),
    .B1(net29),
    .C1(net52),
    .X(_267_));
 sky130_fd_sc_hd__a211o_1 _706_ (.A1(net44),
    .A2(_266_),
    .B1(_267_),
    .C1(net41),
    .X(_268_));
 sky130_fd_sc_hd__a21o_1 _707_ (.A1(_023_),
    .A2(_063_),
    .B1(net21),
    .X(_269_));
 sky130_fd_sc_hd__o22a_1 _708_ (.A1(net26),
    .A2(_050_),
    .B1(_088_),
    .B2(_099_),
    .X(_270_));
 sky130_fd_sc_hd__o311a_1 _709_ (.A1(net22),
    .A2(_054_),
    .A3(_270_),
    .B1(_269_),
    .C1(net37),
    .X(_271_));
 sky130_fd_sc_hd__a21oi_1 _710_ (.A1(_356_),
    .A2(_179_),
    .B1(net21),
    .Y(_272_));
 sky130_fd_sc_hd__nor2_1 _711_ (.A(net37),
    .B(_272_),
    .Y(_273_));
 sky130_fd_sc_hd__o311a_1 _712_ (.A1(_041_),
    .A2(_088_),
    .A3(_099_),
    .B1(_217_),
    .C1(net44),
    .X(_274_));
 sky130_fd_sc_hd__a31o_1 _713_ (.A1(net29),
    .A2(_023_),
    .A3(_063_),
    .B1(net41),
    .X(_275_));
 sky130_fd_sc_hd__o32a_1 _714_ (.A1(net22),
    .A2(_055_),
    .A3(_222_),
    .B1(_274_),
    .B2(_275_),
    .X(_276_));
 sky130_fd_sc_hd__a22o_1 _715_ (.A1(_268_),
    .A2(_271_),
    .B1(_273_),
    .B2(_276_),
    .X(_277_));
 sky130_fd_sc_hd__mux2_1 _716_ (.A0(net25),
    .A1(_249_),
    .S(_277_),
    .X(net17));
 sky130_fd_sc_hd__or2_1 _717_ (.A(_354_),
    .B(_057_),
    .X(_002_));
 sky130_fd_sc_hd__o211a_1 _718_ (.A1(_018_),
    .A2(_022_),
    .B1(net48),
    .C1(_338_),
    .X(_278_));
 sky130_fd_sc_hd__o31ai_1 _719_ (.A1(net48),
    .A2(_354_),
    .A3(_057_),
    .B1(net32),
    .Y(_279_));
 sky130_fd_sc_hd__a21o_1 _720_ (.A1(_351_),
    .A2(_127_),
    .B1(_377_),
    .X(_280_));
 sky130_fd_sc_hd__a31o_1 _721_ (.A1(_341_),
    .A2(_001_),
    .A3(_049_),
    .B1(_239_),
    .X(_281_));
 sky130_fd_sc_hd__o31a_1 _722_ (.A1(_038_),
    .A2(_278_),
    .A3(_279_),
    .B1(net39),
    .X(_282_));
 sky130_fd_sc_hd__nor2_1 _723_ (.A(_057_),
    .B(_179_),
    .Y(_283_));
 sky130_fd_sc_hd__or3_1 _724_ (.A(net60),
    .B(_377_),
    .C(_018_),
    .X(_284_));
 sky130_fd_sc_hd__o311a_1 _725_ (.A1(net22),
    .A2(_062_),
    .A3(_283_),
    .B1(_284_),
    .C1(net34),
    .X(_285_));
 sky130_fd_sc_hd__a31o_1 _726_ (.A1(_280_),
    .A2(_281_),
    .A3(_282_),
    .B1(_285_),
    .X(_286_));
 sky130_fd_sc_hd__a22o_1 _727_ (.A1(net65),
    .A2(_379_),
    .B1(_383_),
    .B2(net56),
    .X(_287_));
 sky130_fd_sc_hd__a211o_1 _728_ (.A1(_101_),
    .A2(_287_),
    .B1(net31),
    .C1(_098_),
    .X(_288_));
 sky130_fd_sc_hd__a31o_1 _729_ (.A1(net57),
    .A2(_089_),
    .A3(_122_),
    .B1(_081_),
    .X(_289_));
 sky130_fd_sc_hd__nand2_1 _730_ (.A(net31),
    .B(_289_),
    .Y(_290_));
 sky130_fd_sc_hd__a21oi_1 _731_ (.A1(_288_),
    .A2(_290_),
    .B1(net20),
    .Y(_291_));
 sky130_fd_sc_hd__nand2_1 _732_ (.A(net36),
    .B(_286_),
    .Y(_292_));
 sky130_fd_sc_hd__o31a_1 _733_ (.A1(_128_),
    .A2(_222_),
    .A3(_235_),
    .B1(_288_),
    .X(_293_));
 sky130_fd_sc_hd__o21a_1 _734_ (.A1(net20),
    .A2(_293_),
    .B1(_286_),
    .X(_294_));
 sky130_fd_sc_hd__o22a_1 _735_ (.A1(_291_),
    .A2(_292_),
    .B1(_294_),
    .B2(net36),
    .X(net3));
 sky130_fd_sc_hd__or3_1 _736_ (.A(net57),
    .B(_360_),
    .C(_021_),
    .X(_295_));
 sky130_fd_sc_hd__a21o_1 _737_ (.A1(_184_),
    .A2(_295_),
    .B1(net21),
    .X(_296_));
 sky130_fd_sc_hd__o32a_1 _738_ (.A1(net27),
    .A2(_345_),
    .A3(_360_),
    .B1(_018_),
    .B2(_022_),
    .X(_297_));
 sky130_fd_sc_hd__or3b_1 _739_ (.A(_342_),
    .B(net22),
    .C_N(_297_),
    .X(_298_));
 sky130_fd_sc_hd__o21a_1 _740_ (.A1(_018_),
    .A2(_055_),
    .B1(_042_),
    .X(_299_));
 sky130_fd_sc_hd__o31a_1 _741_ (.A1(net48),
    .A2(_347_),
    .A3(_023_),
    .B1(net32),
    .X(_300_));
 sky130_fd_sc_hd__o21ai_1 _742_ (.A1(net29),
    .A2(_299_),
    .B1(_300_),
    .Y(_301_));
 sky130_fd_sc_hd__a31oi_1 _743_ (.A1(_296_),
    .A2(_298_),
    .A3(_301_),
    .B1(_328_),
    .Y(_302_));
 sky130_fd_sc_hd__a21oi_1 _744_ (.A1(net28),
    .A2(_002_),
    .B1(_044_),
    .Y(_303_));
 sky130_fd_sc_hd__or4_1 _745_ (.A(_334_),
    .B(net59),
    .C(net68),
    .D(net74),
    .X(_304_));
 sky130_fd_sc_hd__o211a_1 _746_ (.A1(net48),
    .A2(_303_),
    .B1(_304_),
    .C1(_028_),
    .X(_305_));
 sky130_fd_sc_hd__a31o_1 _747_ (.A1(_341_),
    .A2(_349_),
    .A3(_157_),
    .B1(_283_),
    .X(_306_));
 sky130_fd_sc_hd__a22o_1 _748_ (.A1(_148_),
    .A2(_172_),
    .B1(_306_),
    .B2(net46),
    .X(_307_));
 sky130_fd_sc_hd__a211o_1 _749_ (.A1(_029_),
    .A2(_307_),
    .B1(_305_),
    .C1(_302_),
    .X(_308_));
 sky130_fd_sc_hd__mux2_1 _750_ (.A0(_249_),
    .A1(net25),
    .S(_308_),
    .X(net4));
 sky130_fd_sc_hd__mux2_1 _751_ (.A0(_359_),
    .A1(_051_),
    .S(net28),
    .X(_309_));
 sky130_fd_sc_hd__a21o_1 _752_ (.A1(net45),
    .A2(_309_),
    .B1(net42),
    .X(_310_));
 sky130_fd_sc_hd__a211o_1 _753_ (.A1(net28),
    .A2(_051_),
    .B1(_165_),
    .C1(net45),
    .X(_311_));
 sky130_fd_sc_hd__a32o_1 _754_ (.A1(net26),
    .A2(_346_),
    .A3(_018_),
    .B1(_353_),
    .B2(_339_),
    .X(_312_));
 sky130_fd_sc_hd__a21oi_1 _755_ (.A1(_376_),
    .A2(_312_),
    .B1(net34),
    .Y(_313_));
 sky130_fd_sc_hd__and3_1 _756_ (.A(_310_),
    .B(_311_),
    .C(_313_),
    .X(_314_));
 sky130_fd_sc_hd__o21ai_1 _757_ (.A1(_115_),
    .A2(_165_),
    .B1(net29),
    .Y(_315_));
 sky130_fd_sc_hd__o311a_1 _758_ (.A1(net30),
    .A2(_339_),
    .A3(_115_),
    .B1(_315_),
    .C1(_029_),
    .X(_316_));
 sky130_fd_sc_hd__a311o_1 _759_ (.A1(_045_),
    .A2(_078_),
    .A3(_199_),
    .B1(_314_),
    .C1(_316_),
    .X(_317_));
 sky130_fd_sc_hd__a21oi_1 _760_ (.A1(net28),
    .A2(_021_),
    .B1(net25),
    .Y(_318_));
 sky130_fd_sc_hd__mux2_1 _761_ (.A0(net25),
    .A1(_318_),
    .S(_317_),
    .X(net5));
 sky130_fd_sc_hd__or2_1 _762_ (.A(net30),
    .B(_157_),
    .X(_319_));
 sky130_fd_sc_hd__or2_1 _763_ (.A(net45),
    .B(_147_),
    .X(_320_));
 sky130_fd_sc_hd__a221o_1 _764_ (.A1(net33),
    .A2(_046_),
    .B1(_319_),
    .B2(_320_),
    .C1(net34),
    .X(_321_));
 sky130_fd_sc_hd__o21ai_1 _765_ (.A1(_165_),
    .A2(_220_),
    .B1(net30),
    .Y(_322_));
 sky130_fd_sc_hd__a21o_1 _766_ (.A1(_319_),
    .A2(_322_),
    .B1(_030_),
    .X(_323_));
 sky130_fd_sc_hd__o311a_1 _767_ (.A1(net38),
    .A2(_373_),
    .A3(_078_),
    .B1(_321_),
    .C1(_323_),
    .X(_324_));
 sky130_fd_sc_hd__o21a_1 _768_ (.A1(net20),
    .A2(_248_),
    .B1(net25),
    .X(_325_));
 sky130_fd_sc_hd__mux2_1 _769_ (.A0(net35),
    .A1(_325_),
    .S(_324_),
    .X(net6));
 sky130_fd_sc_hd__o211a_1 _770_ (.A1(net45),
    .A2(_147_),
    .B1(net38),
    .C1(net42),
    .X(_326_));
 sky130_fd_sc_hd__a31o_1 _771_ (.A1(_029_),
    .A2(_248_),
    .A3(_319_),
    .B1(_326_),
    .X(_327_));
 sky130_fd_sc_hd__mux2_1 _772_ (.A0(_325_),
    .A1(net35),
    .S(_327_),
    .X(net7));
 sky130_fd_sc_hd__o21a_1 _773_ (.A1(net20),
    .A2(_248_),
    .B1(net35),
    .X(net8));
 sky130_fd_sc_hd__o211ai_1 _774_ (.A1(_347_),
    .A2(_367_),
    .B1(_032_),
    .C1(_338_),
    .Y(_003_));
 sky130_fd_sc_hd__and3_1 _775_ (.A(net50),
    .B(net24),
    .C(_044_),
    .X(_329_));
 sky130_fd_sc_hd__a21o_1 _776_ (.A1(net24),
    .A2(_044_),
    .B1(net49),
    .X(_330_));
 sky130_fd_sc_hd__and2b_1 _777_ (.A_N(_329_),
    .B(_330_),
    .X(_004_));
 sky130_fd_sc_hd__xnor2_1 _778_ (.A(net33),
    .B(_329_),
    .Y(_005_));
 sky130_fd_sc_hd__and3_1 _779_ (.A(net40),
    .B(net43),
    .C(_329_),
    .X(_331_));
 sky130_fd_sc_hd__a21oi_1 _780_ (.A1(net43),
    .A2(_329_),
    .B1(net40),
    .Y(_332_));
 sky130_fd_sc_hd__nor2_1 _781_ (.A(_331_),
    .B(_332_),
    .Y(_006_));
 sky130_fd_sc_hd__xnor2_1 _782_ (.A(net25),
    .B(_331_),
    .Y(_007_));
 sky130_fd_sc_hd__inv_2 _783_ (.A(net1),
    .Y(_009_));
 sky130_fd_sc_hd__inv_2 _784_ (.A(net1),
    .Y(_010_));
 sky130_fd_sc_hd__inv_2 _785_ (.A(net1),
    .Y(_011_));
 sky130_fd_sc_hd__inv_2 _786_ (.A(net1),
    .Y(_012_));
 sky130_fd_sc_hd__inv_2 _787_ (.A(net1),
    .Y(_013_));
 sky130_fd_sc_hd__inv_2 _788_ (.A(net1),
    .Y(_014_));
 sky130_fd_sc_hd__inv_2 _789_ (.A(net1),
    .Y(_015_));
 sky130_fd_sc_hd__dfrtp_1 _790_ (.CLK(clknet_1_0__leaf_clk),
    .D(_000_),
    .RESET_B(_008_),
    .Q(\tcout[0] ));
 sky130_fd_sc_hd__dfrtp_1 _791_ (.CLK(clknet_1_1__leaf_clk),
    .D(net18),
    .RESET_B(_009_),
    .Q(\tcout[1] ));
 sky130_fd_sc_hd__dfrtp_1 _792_ (.CLK(clknet_1_0__leaf_clk),
    .D(_002_),
    .RESET_B(_010_),
    .Q(\tcout[2] ));
 sky130_fd_sc_hd__dfrtp_1 _793_ (.CLK(clknet_1_0__leaf_clk),
    .D(_003_),
    .RESET_B(_011_),
    .Q(\tcout[3] ));
 sky130_fd_sc_hd__dfrtp_1 _794_ (.CLK(clknet_1_0__leaf_clk),
    .D(_004_),
    .RESET_B(_012_),
    .Q(\tcout[4] ));
 sky130_fd_sc_hd__dfrtp_1 _795_ (.CLK(clknet_1_1__leaf_clk),
    .D(_005_),
    .RESET_B(_013_),
    .Q(\tcout[5] ));
 sky130_fd_sc_hd__dfrtp_1 _796_ (.CLK(clknet_1_1__leaf_clk),
    .D(_006_),
    .RESET_B(_014_),
    .Q(\tcout[6] ));
 sky130_fd_sc_hd__dfrtp_1 _797_ (.CLK(clknet_1_1__leaf_clk),
    .D(_007_),
    .RESET_B(_015_),
    .Q(\tcout[7] ));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_160 ();
 sky130_fd_sc_hd__clkbuf_4 input1 (.A(rst),
    .X(net1));
 sky130_fd_sc_hd__buf_2 output2 (.A(net2),
    .X(sine_out[0]));
 sky130_fd_sc_hd__buf_2 output3 (.A(net3),
    .X(sine_out[10]));
 sky130_fd_sc_hd__buf_2 output4 (.A(net4),
    .X(sine_out[11]));
 sky130_fd_sc_hd__buf_2 output5 (.A(net5),
    .X(sine_out[12]));
 sky130_fd_sc_hd__buf_2 output6 (.A(net6),
    .X(sine_out[13]));
 sky130_fd_sc_hd__buf_2 output7 (.A(net7),
    .X(sine_out[14]));
 sky130_fd_sc_hd__buf_2 output8 (.A(net8),
    .X(sine_out[15]));
 sky130_fd_sc_hd__buf_2 output9 (.A(net9),
    .X(sine_out[1]));
 sky130_fd_sc_hd__buf_2 output10 (.A(net10),
    .X(sine_out[2]));
 sky130_fd_sc_hd__buf_2 output11 (.A(net11),
    .X(sine_out[3]));
 sky130_fd_sc_hd__buf_2 output12 (.A(net12),
    .X(sine_out[4]));
 sky130_fd_sc_hd__buf_2 output13 (.A(net13),
    .X(sine_out[5]));
 sky130_fd_sc_hd__buf_2 output14 (.A(net14),
    .X(sine_out[6]));
 sky130_fd_sc_hd__buf_2 output15 (.A(net15),
    .X(sine_out[7]));
 sky130_fd_sc_hd__buf_2 output16 (.A(net16),
    .X(sine_out[8]));
 sky130_fd_sc_hd__buf_2 output17 (.A(net17),
    .X(sine_out[9]));
 sky130_fd_sc_hd__buf_2 fanout18 (.A(_001_),
    .X(net18));
 sky130_fd_sc_hd__buf_1 wire19 (.A(_137_),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_4 fanout20 (.A(_030_),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_4 fanout21 (.A(_377_),
    .X(net21));
 sky130_fd_sc_hd__buf_2 fanout22 (.A(_373_),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_4 fanout23 (.A(_367_),
    .X(net23));
 sky130_fd_sc_hd__buf_2 fanout24 (.A(_352_),
    .X(net24));
 sky130_fd_sc_hd__buf_2 fanout25 (.A(_337_),
    .X(net25));
 sky130_fd_sc_hd__buf_2 fanout26 (.A(net28),
    .X(net26));
 sky130_fd_sc_hd__buf_2 fanout27 (.A(net28),
    .X(net27));
 sky130_fd_sc_hd__buf_2 fanout28 (.A(_335_),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_4 fanout29 (.A(net31),
    .X(net29));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout30 (.A(net31),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_4 fanout31 (.A(_334_),
    .X(net31));
 sky130_fd_sc_hd__buf_4 fanout32 (.A(_333_),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_2 fanout33 (.A(_333_),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_4 fanout34 (.A(_328_),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_4 fanout35 (.A(\tcout[7] ),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_2 fanout36 (.A(\tcout[7] ),
    .X(net36));
 sky130_fd_sc_hd__buf_2 fanout37 (.A(net40),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_2 fanout38 (.A(net40),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_4 fanout39 (.A(net40),
    .X(net39));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout40 (.A(\tcout[6] ),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_4 fanout41 (.A(net43),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_2 fanout42 (.A(net43),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_4 fanout43 (.A(\tcout[5] ),
    .X(net43));
 sky130_fd_sc_hd__buf_2 fanout44 (.A(net47),
    .X(net44));
 sky130_fd_sc_hd__buf_2 fanout45 (.A(net47),
    .X(net45));
 sky130_fd_sc_hd__buf_2 fanout46 (.A(net47),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_2 fanout47 (.A(\tcout[4] ),
    .X(net47));
 sky130_fd_sc_hd__buf_2 fanout48 (.A(net50),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_4 fanout49 (.A(net50),
    .X(net49));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout50 (.A(\tcout[4] ),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_4 fanout51 (.A(net55),
    .X(net51));
 sky130_fd_sc_hd__buf_2 fanout52 (.A(net54),
    .X(net52));
 sky130_fd_sc_hd__buf_1 fanout53 (.A(net54),
    .X(net53));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout54 (.A(net55),
    .X(net54));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout55 (.A(net60),
    .X(net55));
 sky130_fd_sc_hd__buf_2 fanout56 (.A(net57),
    .X(net56));
 sky130_fd_sc_hd__buf_2 fanout57 (.A(net60),
    .X(net57));
 sky130_fd_sc_hd__buf_2 fanout58 (.A(net60),
    .X(net58));
 sky130_fd_sc_hd__buf_1 fanout59 (.A(net60),
    .X(net59));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout60 (.A(\tcout[3] ),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_8 fanout61 (.A(net62),
    .X(net61));
 sky130_fd_sc_hd__buf_2 fanout62 (.A(net69),
    .X(net62));
 sky130_fd_sc_hd__buf_2 fanout63 (.A(net64),
    .X(net63));
 sky130_fd_sc_hd__buf_2 fanout64 (.A(net69),
    .X(net64));
 sky130_fd_sc_hd__buf_2 fanout65 (.A(net68),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_2 fanout66 (.A(net68),
    .X(net66));
 sky130_fd_sc_hd__buf_2 fanout67 (.A(net68),
    .X(net67));
 sky130_fd_sc_hd__buf_1 fanout68 (.A(net69),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_2 fanout69 (.A(\tcout[2] ),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_8 fanout70 (.A(net72),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_4 fanout71 (.A(net72),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_2 fanout72 (.A(\tcout[1] ),
    .X(net72));
 sky130_fd_sc_hd__buf_2 fanout73 (.A(net74),
    .X(net73));
 sky130_fd_sc_hd__buf_2 fanout74 (.A(\tcout[1] ),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_8 fanout75 (.A(net76),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_4 fanout76 (.A(net79),
    .X(net76));
 sky130_fd_sc_hd__buf_2 fanout77 (.A(net79),
    .X(net77));
 sky130_fd_sc_hd__buf_2 fanout78 (.A(net79),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_2 fanout79 (.A(\tcout[0] ),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .X(clknet_1_1__leaf_clk));
 sky130_ef_sc_hd__decap_12 FILLER_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_140 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_140 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_18 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_185 ();
endmodule
