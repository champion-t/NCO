VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO counter
  CLASS BLOCK ;
  FOREIGN counter ;
  ORIGIN 0.000 0.000 ;
  SIZE 560.000 BY 370.000 ;
  PIN addr0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END addr0[0]
  PIN addr0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 4.000 ;
    END
  END addr0[1]
  PIN addr0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END addr0[2]
  PIN addr0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END addr0[3]
  PIN addr0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END addr0[4]
  PIN addr0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 4.000 191.040 ;
    END
  END addr0[5]
  PIN addr0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.240 4.000 197.840 ;
    END
  END addr0[6]
  PIN addr0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 207.440 4.000 208.040 ;
    END
  END addr0[7]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 556.000 51.040 560.000 51.640 ;
    END
  END clk
  PIN csb0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END csb0
  PIN din0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END din0[0]
  PIN din0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met2 ;
        RECT 186.850 0.000 187.130 4.000 ;
    END
  END din0[10]
  PIN din0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END din0[11]
  PIN din0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met2 ;
        RECT 199.730 0.000 200.010 4.000 ;
    END
  END din0[12]
  PIN din0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met2 ;
        RECT 206.170 0.000 206.450 4.000 ;
    END
  END din0[13]
  PIN din0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met2 ;
        RECT 209.390 0.000 209.670 4.000 ;
    END
  END din0[14]
  PIN din0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met2 ;
        RECT 215.830 0.000 216.110 4.000 ;
    END
  END din0[15]
  PIN din0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END din0[1]
  PIN din0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met2 ;
        RECT 141.770 0.000 142.050 4.000 ;
    END
  END din0[2]
  PIN din0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 4.000 ;
    END
  END din0[3]
  PIN din0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met2 ;
        RECT 151.430 0.000 151.710 4.000 ;
    END
  END din0[4]
  PIN din0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met2 ;
        RECT 157.870 0.000 158.150 4.000 ;
    END
  END din0[5]
  PIN din0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END din0[6]
  PIN din0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 4.000 ;
    END
  END din0[7]
  PIN din0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END din0[8]
  PIN din0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.600000 ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 4.000 ;
    END
  END din0[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 556.000 156.440 560.000 157.040 ;
    END
  END rst
  PIN sine_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 222.270 366.000 222.550 370.000 ;
    END
  END sine_out[0]
  PIN sine_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 328.530 366.000 328.810 370.000 ;
    END
  END sine_out[10]
  PIN sine_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 338.190 366.000 338.470 370.000 ;
    END
  END sine_out[11]
  PIN sine_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 347.850 366.000 348.130 370.000 ;
    END
  END sine_out[12]
  PIN sine_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 357.510 366.000 357.790 370.000 ;
    END
  END sine_out[13]
  PIN sine_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 370.390 366.000 370.670 370.000 ;
    END
  END sine_out[14]
  PIN sine_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 386.490 366.000 386.770 370.000 ;
    END
  END sine_out[15]
  PIN sine_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 235.150 366.000 235.430 370.000 ;
    END
  END sine_out[1]
  PIN sine_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 248.030 366.000 248.310 370.000 ;
    END
  END sine_out[2]
  PIN sine_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 257.690 366.000 257.970 370.000 ;
    END
  END sine_out[3]
  PIN sine_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 267.350 366.000 267.630 370.000 ;
    END
  END sine_out[4]
  PIN sine_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 277.010 366.000 277.290 370.000 ;
    END
  END sine_out[5]
  PIN sine_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 286.670 366.000 286.950 370.000 ;
    END
  END sine_out[6]
  PIN sine_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 296.330 366.000 296.610 370.000 ;
    END
  END sine_out[7]
  PIN sine_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 305.990 366.000 306.270 370.000 ;
    END
  END sine_out[8]
  PIN sine_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 315.650 366.000 315.930 370.000 ;
    END
  END sine_out[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 359.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 39.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 328.250 176.240 359.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 40.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 328.880 329.840 359.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 40.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 328.250 483.440 359.280 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 26.730 554.540 28.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 179.910 554.540 181.510 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 333.090 554.540 334.690 ;
    END
    PORT
      LAYER met4 ;
        RECT 535.100 35.120 536.700 332.080 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 359.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 10.640 179.540 40.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 328.250 179.540 359.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 331.540 10.640 333.140 40.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 331.540 328.250 333.140 359.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 485.140 10.640 486.740 40.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 485.140 328.250 486.740 359.280 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 30.030 554.540 31.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 183.210 554.540 184.810 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 336.390 554.540 337.990 ;
    END
    PORT
      LAYER met4 ;
        RECT 538.780 35.120 540.380 332.080 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 554.490 359.125 ;
      LAYER li1 ;
        RECT 5.520 10.795 554.300 359.125 ;
      LAYER met1 ;
        RECT 5.520 10.640 554.300 359.280 ;
      LAYER met2 ;
        RECT 21.070 365.720 221.990 366.000 ;
        RECT 222.830 365.720 234.870 366.000 ;
        RECT 235.710 365.720 247.750 366.000 ;
        RECT 248.590 365.720 257.410 366.000 ;
        RECT 258.250 365.720 267.070 366.000 ;
        RECT 267.910 365.720 276.730 366.000 ;
        RECT 277.570 365.720 286.390 366.000 ;
        RECT 287.230 365.720 296.050 366.000 ;
        RECT 296.890 365.720 305.710 366.000 ;
        RECT 306.550 365.720 315.370 366.000 ;
        RECT 316.210 365.720 328.250 366.000 ;
        RECT 329.090 365.720 337.910 366.000 ;
        RECT 338.750 365.720 347.570 366.000 ;
        RECT 348.410 365.720 357.230 366.000 ;
        RECT 358.070 365.720 370.110 366.000 ;
        RECT 370.950 365.720 386.210 366.000 ;
        RECT 387.050 365.720 552.830 366.000 ;
        RECT 21.070 4.280 552.830 365.720 ;
        RECT 21.070 4.000 115.730 4.280 ;
        RECT 116.570 4.000 122.170 4.280 ;
        RECT 123.010 4.000 128.610 4.280 ;
        RECT 129.450 4.000 135.050 4.280 ;
        RECT 135.890 4.000 141.490 4.280 ;
        RECT 142.330 4.000 144.710 4.280 ;
        RECT 145.550 4.000 151.150 4.280 ;
        RECT 151.990 4.000 157.590 4.280 ;
        RECT 158.430 4.000 164.030 4.280 ;
        RECT 164.870 4.000 170.470 4.280 ;
        RECT 171.310 4.000 176.910 4.280 ;
        RECT 177.750 4.000 180.130 4.280 ;
        RECT 180.970 4.000 186.570 4.280 ;
        RECT 187.410 4.000 193.010 4.280 ;
        RECT 193.850 4.000 199.450 4.280 ;
        RECT 200.290 4.000 205.890 4.280 ;
        RECT 206.730 4.000 209.110 4.280 ;
        RECT 209.950 4.000 215.550 4.280 ;
        RECT 216.390 4.000 552.830 4.280 ;
      LAYER met3 ;
        RECT 4.000 208.440 556.000 359.205 ;
        RECT 4.400 207.040 556.000 208.440 ;
        RECT 4.000 198.240 556.000 207.040 ;
        RECT 4.400 196.840 556.000 198.240 ;
        RECT 4.000 191.440 556.000 196.840 ;
        RECT 4.400 190.040 556.000 191.440 ;
        RECT 4.000 184.640 556.000 190.040 ;
        RECT 4.400 183.240 556.000 184.640 ;
        RECT 4.000 177.840 556.000 183.240 ;
        RECT 4.400 176.440 556.000 177.840 ;
        RECT 4.000 171.040 556.000 176.440 ;
        RECT 4.400 169.640 556.000 171.040 ;
        RECT 4.000 157.440 556.000 169.640 ;
        RECT 4.000 156.040 555.600 157.440 ;
        RECT 4.000 79.240 556.000 156.040 ;
        RECT 4.400 77.840 556.000 79.240 ;
        RECT 4.000 52.040 556.000 77.840 ;
        RECT 4.000 50.640 555.600 52.040 ;
        RECT 4.000 6.295 556.000 50.640 ;
      LAYER met4 ;
        RECT 50.000 327.850 174.240 335.745 ;
        RECT 176.640 327.850 177.540 335.745 ;
        RECT 179.940 328.480 327.840 335.745 ;
        RECT 330.240 328.480 331.140 335.745 ;
        RECT 179.940 327.850 331.140 328.480 ;
        RECT 333.540 327.850 481.440 335.745 ;
        RECT 483.840 327.850 484.740 335.745 ;
        RECT 487.140 327.850 509.900 335.745 ;
        RECT 50.000 40.720 509.900 327.850 ;
        RECT 50.000 39.800 177.540 40.720 ;
        RECT 50.000 10.240 174.240 39.800 ;
        RECT 176.640 10.240 177.540 39.800 ;
        RECT 179.940 10.240 327.840 40.720 ;
        RECT 330.240 10.240 331.140 40.720 ;
        RECT 333.540 10.240 481.440 40.720 ;
        RECT 483.840 10.240 484.740 40.720 ;
        RECT 487.140 10.240 509.900 40.720 ;
        RECT 50.000 6.295 509.900 10.240 ;
  END
END counter
END LIBRARY

