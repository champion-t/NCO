module counter (clk,
    rst,
    sine_out,
    VPWR,
    VGND);
 input clk;
 input rst;
 output [15:0] sine_out;
 inout VPWR;
 inout VGND;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire _369_;
 wire _370_;
 wire _371_;
 wire _372_;
 wire _373_;
 wire _374_;
 wire _375_;
 wire _376_;
 wire _377_;
 wire _378_;
 wire _379_;
 wire _380_;
 wire _381_;
 wire _382_;
 wire _383_;
 wire _384_;
 wire _385_;
 wire _386_;
 wire \tcout[0] ;
 wire \tcout[1] ;
 wire \tcout[2] ;
 wire \tcout[3] ;
 wire \tcout[4] ;
 wire \tcout[5] ;
 wire \tcout[6] ;
 wire \tcout[7] ;

 sky130_fd_sc_hd__inv_2 _387_ (.A(\tcout[0] ),
    .Y(_000_));
 sky130_fd_sc_hd__inv_2 _388_ (.A(\tcout[6] ),
    .Y(_328_));
 sky130_fd_sc_hd__inv_2 _389_ (.A(\tcout[5] ),
    .Y(_333_));
 sky130_fd_sc_hd__inv_2 _390_ (.A(\tcout[4] ),
    .Y(_334_));
 sky130_fd_sc_hd__inv_2 _391_ (.A(\tcout[3] ),
    .Y(_335_));
 sky130_fd_sc_hd__inv_2 _392_ (.A(\tcout[2] ),
    .Y(_336_));
 sky130_fd_sc_hd__inv_2 _393_ (.A(\tcout[7] ),
    .Y(_337_));
 sky130_fd_sc_hd__inv_2 _394_ (.A(rst),
    .Y(_008_));
 sky130_fd_sc_hd__nand2b_2 _395_ (.A_N(\tcout[1] ),
    .B(\tcout[3] ),
    .Y(_338_));
 sky130_fd_sc_hd__and2b_2 _396_ (.A_N(\tcout[2] ),
    .B(\tcout[3] ),
    .X(_339_));
 sky130_fd_sc_hd__nor2_2 _397_ (.A(\tcout[2] ),
    .B(\tcout[1] ),
    .Y(_340_));
 sky130_fd_sc_hd__or2_2 _398_ (.A(\tcout[2] ),
    .B(\tcout[1] ),
    .X(_341_));
 sky130_fd_sc_hd__nor3b_2 _399_ (.A(\tcout[2] ),
    .B(\tcout[1] ),
    .C_N(\tcout[3] ),
    .Y(_342_));
 sky130_fd_sc_hd__nand2_2 _400_ (.A(\tcout[3] ),
    .B(_340_),
    .Y(_343_));
 sky130_fd_sc_hd__and2b_2 _401_ (.A_N(\tcout[0] ),
    .B(\tcout[2] ),
    .X(_344_));
 sky130_fd_sc_hd__and2b_2 _402_ (.A_N(\tcout[2] ),
    .B(\tcout[0] ),
    .X(_345_));
 sky130_fd_sc_hd__nand2b_2 _403_ (.A_N(\tcout[2] ),
    .B(\tcout[0] ),
    .Y(_346_));
 sky130_fd_sc_hd__nand2_2 _404_ (.A(\tcout[0] ),
    .B(\tcout[2] ),
    .Y(_347_));
 sky130_fd_sc_hd__nor2_2 _405_ (.A(\tcout[0] ),
    .B(\tcout[2] ),
    .Y(_348_));
 sky130_fd_sc_hd__or2_2 _406_ (.A(\tcout[0] ),
    .B(\tcout[2] ),
    .X(_349_));
 sky130_fd_sc_hd__xnor2_2 _407_ (.A(\tcout[0] ),
    .B(\tcout[2] ),
    .Y(_350_));
 sky130_fd_sc_hd__nand2_2 _408_ (.A(\tcout[3] ),
    .B(_350_),
    .Y(_351_));
 sky130_fd_sc_hd__and2_2 _409_ (.A(\tcout[0] ),
    .B(\tcout[1] ),
    .X(_352_));
 sky130_fd_sc_hd__nand2_2 _410_ (.A(\tcout[0] ),
    .B(\tcout[1] ),
    .Y(_353_));
 sky130_fd_sc_hd__and3b_2 _411_ (.A_N(\tcout[2] ),
    .B(\tcout[1] ),
    .C(\tcout[0] ),
    .X(_354_));
 sky130_fd_sc_hd__a211o_2 _412_ (.A1(\tcout[3] ),
    .A2(_350_),
    .B1(_342_),
    .C1(\tcout[4] ),
    .X(_355_));
 sky130_fd_sc_hd__or2_2 _413_ (.A(\tcout[3] ),
    .B(\tcout[1] ),
    .X(_356_));
 sky130_fd_sc_hd__nand2_2 _414_ (.A(_335_),
    .B(\tcout[2] ),
    .Y(_357_));
 sky130_fd_sc_hd__a21oi_2 _415_ (.A1(\tcout[1] ),
    .A2(_347_),
    .B1(\tcout[3] ),
    .Y(_358_));
 sky130_fd_sc_hd__nand2_2 _416_ (.A(\tcout[2] ),
    .B(\tcout[1] ),
    .Y(_359_));
 sky130_fd_sc_hd__and2b_2 _417_ (.A_N(\tcout[1] ),
    .B(\tcout[2] ),
    .X(_360_));
 sky130_fd_sc_hd__nand2b_2 _418_ (.A_N(\tcout[1] ),
    .B(\tcout[2] ),
    .Y(_361_));
 sky130_fd_sc_hd__nand2_2 _419_ (.A(_335_),
    .B(_360_),
    .Y(_362_));
 sky130_fd_sc_hd__nand2_2 _420_ (.A(_346_),
    .B(_362_),
    .Y(_363_));
 sky130_fd_sc_hd__a2bb2o_2 _421_ (.A1_N(_355_),
    .A2_N(_358_),
    .B1(_363_),
    .B2(\tcout[4] ),
    .X(_364_));
 sky130_fd_sc_hd__nand2_2 _422_ (.A(\tcout[2] ),
    .B(_352_),
    .Y(_365_));
 sky130_fd_sc_hd__and2b_2 _423_ (.A_N(\tcout[3] ),
    .B(\tcout[1] ),
    .X(_366_));
 sky130_fd_sc_hd__nand2b_2 _424_ (.A_N(\tcout[3] ),
    .B(\tcout[1] ),
    .Y(_367_));
 sky130_fd_sc_hd__o21bai_2 _425_ (.A1(\tcout[2] ),
    .A2(\tcout[1] ),
    .B1_N(\tcout[3] ),
    .Y(_368_));
 sky130_fd_sc_hd__a21o_2 _426_ (.A1(\tcout[2] ),
    .A2(_352_),
    .B1(_368_),
    .X(_369_));
 sky130_fd_sc_hd__nand2_2 _427_ (.A(\tcout[0] ),
    .B(\tcout[3] ),
    .Y(_370_));
 sky130_fd_sc_hd__nand2_2 _428_ (.A(\tcout[3] ),
    .B(_352_),
    .Y(_371_));
 sky130_fd_sc_hd__nor2_2 _429_ (.A(_333_),
    .B(\tcout[4] ),
    .Y(_372_));
 sky130_fd_sc_hd__nand2b_2 _430_ (.A_N(\tcout[4] ),
    .B(\tcout[5] ),
    .Y(_373_));
 sky130_fd_sc_hd__or2_2 _431_ (.A(\tcout[0] ),
    .B(\tcout[1] ),
    .X(_374_));
 sky130_fd_sc_hd__xnor2_2 _432_ (.A(\tcout[0] ),
    .B(\tcout[1] ),
    .Y(_375_));
 sky130_fd_sc_hd__inv_2 _433_ (.A(_375_),
    .Y(_001_));
 sky130_fd_sc_hd__nor2_2 _434_ (.A(_333_),
    .B(_334_),
    .Y(_376_));
 sky130_fd_sc_hd__nand2_2 _435_ (.A(\tcout[5] ),
    .B(\tcout[4] ),
    .Y(_377_));
 sky130_fd_sc_hd__and2b_2 _436_ (.A_N(\tcout[0] ),
    .B(\tcout[1] ),
    .X(_378_));
 sky130_fd_sc_hd__nand2b_2 _437_ (.A_N(\tcout[0] ),
    .B(\tcout[1] ),
    .Y(_379_));
 sky130_fd_sc_hd__and2b_2 _438_ (.A_N(\tcout[2] ),
    .B(\tcout[1] ),
    .X(_380_));
 sky130_fd_sc_hd__nand2b_2 _439_ (.A_N(\tcout[2] ),
    .B(\tcout[1] ),
    .Y(_381_));
 sky130_fd_sc_hd__and2b_2 _440_ (.A_N(\tcout[1] ),
    .B(\tcout[0] ),
    .X(_382_));
 sky130_fd_sc_hd__nand2b_2 _441_ (.A_N(\tcout[1] ),
    .B(\tcout[0] ),
    .Y(_383_));
 sky130_fd_sc_hd__nand2_2 _442_ (.A(_339_),
    .B(_375_),
    .Y(_384_));
 sky130_fd_sc_hd__o311a_2 _443_ (.A1(\tcout[3] ),
    .A2(_344_),
    .A3(_354_),
    .B1(_384_),
    .C1(\tcout[4] ),
    .X(_385_));
 sky130_fd_sc_hd__a31o_2 _444_ (.A1(_334_),
    .A2(_369_),
    .A3(_371_),
    .B1(_385_),
    .X(_386_));
 sky130_fd_sc_hd__mux2_1 _445_ (.A0(_364_),
    .A1(_386_),
    .S(\tcout[5] ),
    .X(_016_));
 sky130_fd_sc_hd__a21o_2 _446_ (.A1(_341_),
    .A2(_001_),
    .B1(_335_),
    .X(_017_));
 sky130_fd_sc_hd__xnor2_2 _447_ (.A(\tcout[2] ),
    .B(\tcout[1] ),
    .Y(_018_));
 sky130_fd_sc_hd__nor2_2 _448_ (.A(_345_),
    .B(_018_),
    .Y(_019_));
 sky130_fd_sc_hd__o211ai_2 _449_ (.A1(\tcout[3] ),
    .A2(_019_),
    .B1(_017_),
    .C1(\tcout[4] ),
    .Y(_020_));
 sky130_fd_sc_hd__nor3_2 _450_ (.A(\tcout[0] ),
    .B(\tcout[2] ),
    .C(\tcout[1] ),
    .Y(_021_));
 sky130_fd_sc_hd__a21o_2 _451_ (.A1(\tcout[0] ),
    .A2(\tcout[2] ),
    .B1(\tcout[3] ),
    .X(_022_));
 sky130_fd_sc_hd__nand2_2 _452_ (.A(\tcout[3] ),
    .B(\tcout[1] ),
    .Y(_023_));
 sky130_fd_sc_hd__nand2_2 _453_ (.A(\tcout[3] ),
    .B(_378_),
    .Y(_024_));
 sky130_fd_sc_hd__and3_2 _454_ (.A(\tcout[3] ),
    .B(_353_),
    .C(_361_),
    .X(_025_));
 sky130_fd_sc_hd__nor2_2 _455_ (.A(\tcout[4] ),
    .B(_025_),
    .Y(_026_));
 sky130_fd_sc_hd__o21ai_2 _456_ (.A1(_021_),
    .A2(_022_),
    .B1(_026_),
    .Y(_027_));
 sky130_fd_sc_hd__nor2_2 _457_ (.A(\tcout[6] ),
    .B(_333_),
    .Y(_028_));
 sky130_fd_sc_hd__nor2_2 _458_ (.A(\tcout[6] ),
    .B(\tcout[5] ),
    .Y(_029_));
 sky130_fd_sc_hd__or2_2 _459_ (.A(\tcout[6] ),
    .B(\tcout[5] ),
    .X(_030_));
 sky130_fd_sc_hd__a21boi_2 _460_ (.A1(\tcout[0] ),
    .A2(\tcout[2] ),
    .B1_N(\tcout[3] ),
    .Y(_031_));
 sky130_fd_sc_hd__a21bo_2 _461_ (.A1(\tcout[0] ),
    .A2(\tcout[2] ),
    .B1_N(\tcout[3] ),
    .X(_032_));
 sky130_fd_sc_hd__o311a_2 _462_ (.A1(_340_),
    .A2(_382_),
    .A3(_031_),
    .B1(_343_),
    .C1(\tcout[4] ),
    .X(_033_));
 sky130_fd_sc_hd__nand2_2 _463_ (.A(\tcout[3] ),
    .B(_019_),
    .Y(_034_));
 sky130_fd_sc_hd__and3b_2 _464_ (.A_N(\tcout[1] ),
    .B(\tcout[2] ),
    .C(\tcout[0] ),
    .X(_035_));
 sky130_fd_sc_hd__nand3b_2 _465_ (.A_N(\tcout[1] ),
    .B(\tcout[2] ),
    .C(\tcout[0] ),
    .Y(_036_));
 sky130_fd_sc_hd__nand2_2 _466_ (.A(_335_),
    .B(_036_),
    .Y(_037_));
 sky130_fd_sc_hd__nor2_2 _467_ (.A(\tcout[4] ),
    .B(\tcout[3] ),
    .Y(_038_));
 sky130_fd_sc_hd__a31o_2 _468_ (.A1(_334_),
    .A2(_034_),
    .A3(_037_),
    .B1(_033_),
    .X(_039_));
 sky130_fd_sc_hd__a32o_2 _469_ (.A1(_020_),
    .A2(_027_),
    .A3(_028_),
    .B1(_029_),
    .B2(_039_),
    .X(_040_));
 sky130_fd_sc_hd__o21bai_2 _470_ (.A1(_328_),
    .A2(_016_),
    .B1_N(_040_),
    .Y(sine_out[0]));
 sky130_fd_sc_hd__nor2_2 _471_ (.A(\tcout[3] ),
    .B(\tcout[2] ),
    .Y(_041_));
 sky130_fd_sc_hd__or2_2 _472_ (.A(\tcout[3] ),
    .B(\tcout[2] ),
    .X(_042_));
 sky130_fd_sc_hd__a221o_2 _473_ (.A1(_018_),
    .A2(_031_),
    .B1(_041_),
    .B2(_352_),
    .C1(_334_),
    .X(_043_));
 sky130_fd_sc_hd__and2_2 _474_ (.A(\tcout[3] ),
    .B(\tcout[2] ),
    .X(_044_));
 sky130_fd_sc_hd__nand2_2 _475_ (.A(\tcout[3] ),
    .B(\tcout[2] ),
    .Y(_045_));
 sky130_fd_sc_hd__nand2_2 _476_ (.A(\tcout[1] ),
    .B(_044_),
    .Y(_046_));
 sky130_fd_sc_hd__a32oi_2 _477_ (.A1(\tcout[0] ),
    .A2(_341_),
    .A3(_046_),
    .B1(_031_),
    .B2(_001_),
    .Y(_047_));
 sky130_fd_sc_hd__o21ai_2 _478_ (.A1(\tcout[4] ),
    .A2(_047_),
    .B1(_043_),
    .Y(_048_));
 sky130_fd_sc_hd__nand2_2 _479_ (.A(\tcout[3] ),
    .B(_359_),
    .Y(_049_));
 sky130_fd_sc_hd__o21ai_2 _480_ (.A1(\tcout[0] ),
    .A2(\tcout[1] ),
    .B1(\tcout[2] ),
    .Y(_050_));
 sky130_fd_sc_hd__o21a_2 _481_ (.A1(\tcout[0] ),
    .A2(\tcout[1] ),
    .B1(\tcout[2] ),
    .X(_051_));
 sky130_fd_sc_hd__o21ai_2 _482_ (.A1(\tcout[0] ),
    .A2(\tcout[2] ),
    .B1(\tcout[3] ),
    .Y(_052_));
 sky130_fd_sc_hd__a2bb2o_2 _483_ (.A1_N(_051_),
    .A2_N(_052_),
    .B1(_335_),
    .B2(_361_),
    .X(_053_));
 sky130_fd_sc_hd__nor2_2 _484_ (.A(_383_),
    .B(_045_),
    .Y(_054_));
 sky130_fd_sc_hd__and2b_2 _485_ (.A_N(\tcout[3] ),
    .B(\tcout[0] ),
    .X(_055_));
 sky130_fd_sc_hd__nand2_2 _486_ (.A(\tcout[2] ),
    .B(_353_),
    .Y(_056_));
 sky130_fd_sc_hd__a21boi_2 _487_ (.A1(\tcout[0] ),
    .A2(\tcout[1] ),
    .B1_N(\tcout[2] ),
    .Y(_057_));
 sky130_fd_sc_hd__a31o_2 _488_ (.A1(\tcout[0] ),
    .A2(_335_),
    .A3(_018_),
    .B1(_054_),
    .X(_058_));
 sky130_fd_sc_hd__a221o_2 _489_ (.A1(_372_),
    .A2(_053_),
    .B1(_058_),
    .B2(_376_),
    .C1(\tcout[6] ),
    .X(_059_));
 sky130_fd_sc_hd__a21o_2 _490_ (.A1(_333_),
    .A2(_048_),
    .B1(_059_),
    .X(_060_));
 sky130_fd_sc_hd__a21o_2 _491_ (.A1(\tcout[0] ),
    .A2(_018_),
    .B1(_335_),
    .X(_061_));
 sky130_fd_sc_hd__nor2_2 _492_ (.A(\tcout[3] ),
    .B(_375_),
    .Y(_062_));
 sky130_fd_sc_hd__nand2_2 _493_ (.A(_335_),
    .B(_001_),
    .Y(_063_));
 sky130_fd_sc_hd__a31o_2 _494_ (.A1(_357_),
    .A2(_061_),
    .A3(_063_),
    .B1(\tcout[4] ),
    .X(_064_));
 sky130_fd_sc_hd__nand2_2 _495_ (.A(\tcout[2] ),
    .B(_379_),
    .Y(_065_));
 sky130_fd_sc_hd__o31a_2 _496_ (.A1(\tcout[3] ),
    .A2(_336_),
    .A3(_378_),
    .B1(\tcout[4] ),
    .X(_066_));
 sky130_fd_sc_hd__nand2_2 _497_ (.A(\tcout[3] ),
    .B(_374_),
    .Y(_067_));
 sky130_fd_sc_hd__o21ai_2 _498_ (.A1(_354_),
    .A2(_067_),
    .B1(_066_),
    .Y(_068_));
 sky130_fd_sc_hd__and3_2 _499_ (.A(_333_),
    .B(_064_),
    .C(_068_),
    .X(_069_));
 sky130_fd_sc_hd__o32a_2 _500_ (.A1(_335_),
    .A2(_345_),
    .A3(_382_),
    .B1(_356_),
    .B2(_350_),
    .X(_070_));
 sky130_fd_sc_hd__a21bo_2 _501_ (.A1(_338_),
    .A2(_367_),
    .B1_N(_350_),
    .X(_071_));
 sky130_fd_sc_hd__a221o_2 _502_ (.A1(_376_),
    .A2(_070_),
    .B1(_071_),
    .B2(_372_),
    .C1(_328_),
    .X(_072_));
 sky130_fd_sc_hd__o21a_2 _503_ (.A1(_069_),
    .A2(_072_),
    .B1(_337_),
    .X(_073_));
 sky130_fd_sc_hd__a221o_2 _504_ (.A1(\tcout[3] ),
    .A2(\tcout[1] ),
    .B1(_361_),
    .B2(_055_),
    .C1(_054_),
    .X(_074_));
 sky130_fd_sc_hd__a21o_2 _505_ (.A1(_347_),
    .A2(_349_),
    .B1(_049_),
    .X(_075_));
 sky130_fd_sc_hd__nor2_2 _506_ (.A(\tcout[4] ),
    .B(_055_),
    .Y(_076_));
 sky130_fd_sc_hd__a32o_2 _507_ (.A1(_362_),
    .A2(_075_),
    .A3(_076_),
    .B1(_074_),
    .B2(\tcout[4] ),
    .X(_077_));
 sky130_fd_sc_hd__a211o_2 _508_ (.A1(\tcout[0] ),
    .A2(\tcout[1] ),
    .B1(\tcout[2] ),
    .C1(\tcout[3] ),
    .X(_078_));
 sky130_fd_sc_hd__a21o_2 _509_ (.A1(_336_),
    .A2(_375_),
    .B1(_032_),
    .X(_079_));
 sky130_fd_sc_hd__a21o_2 _510_ (.A1(_078_),
    .A2(_079_),
    .B1(_373_),
    .X(_080_));
 sky130_fd_sc_hd__a21oi_2 _511_ (.A1(_367_),
    .A2(_042_),
    .B1(_350_),
    .Y(_081_));
 sky130_fd_sc_hd__o21ba_2 _512_ (.A1(_338_),
    .A2(_344_),
    .B1_N(_081_),
    .X(_082_));
 sky130_fd_sc_hd__o211a_2 _513_ (.A1(_377_),
    .A2(_082_),
    .B1(_080_),
    .C1(\tcout[6] ),
    .X(_083_));
 sky130_fd_sc_hd__o21ai_2 _514_ (.A1(\tcout[5] ),
    .A2(_077_),
    .B1(_083_),
    .Y(_084_));
 sky130_fd_sc_hd__o211ai_2 _515_ (.A1(\tcout[3] ),
    .A2(_353_),
    .B1(_351_),
    .C1(_334_),
    .Y(_085_));
 sky130_fd_sc_hd__or2_2 _516_ (.A(\tcout[0] ),
    .B(_368_),
    .X(_086_));
 sky130_fd_sc_hd__a31oi_2 _517_ (.A1(\tcout[4] ),
    .A2(_359_),
    .A3(_086_),
    .B1(\tcout[5] ),
    .Y(_087_));
 sky130_fd_sc_hd__nor2_2 _518_ (.A(\tcout[2] ),
    .B(_375_),
    .Y(_088_));
 sky130_fd_sc_hd__nand2_2 _519_ (.A(_336_),
    .B(_001_),
    .Y(_089_));
 sky130_fd_sc_hd__a21o_2 _520_ (.A1(_065_),
    .A2(_089_),
    .B1(\tcout[3] ),
    .X(_090_));
 sky130_fd_sc_hd__nor2_2 _521_ (.A(_347_),
    .B(_367_),
    .Y(_091_));
 sky130_fd_sc_hd__a31o_2 _522_ (.A1(_347_),
    .A2(_367_),
    .A3(_383_),
    .B1(_091_),
    .X(_092_));
 sky130_fd_sc_hd__a221o_2 _523_ (.A1(_085_),
    .A2(_087_),
    .B1(_092_),
    .B2(_372_),
    .C1(\tcout[6] ),
    .X(_093_));
 sky130_fd_sc_hd__a31o_2 _524_ (.A1(_376_),
    .A2(_024_),
    .A3(_090_),
    .B1(_093_),
    .X(_094_));
 sky130_fd_sc_hd__a32o_2 _525_ (.A1(\tcout[7] ),
    .A2(_084_),
    .A3(_094_),
    .B1(_060_),
    .B2(_073_),
    .X(sine_out[1]));
 sky130_fd_sc_hd__o21ai_2 _526_ (.A1(\tcout[2] ),
    .A2(\tcout[1] ),
    .B1(\tcout[3] ),
    .Y(_095_));
 sky130_fd_sc_hd__a21oi_2 _527_ (.A1(\tcout[2] ),
    .A2(_001_),
    .B1(_095_),
    .Y(_096_));
 sky130_fd_sc_hd__a211oi_2 _528_ (.A1(_341_),
    .A2(_062_),
    .B1(_096_),
    .C1(_373_),
    .Y(_097_));
 sky130_fd_sc_hd__nor3b_2 _529_ (.A(\tcout[0] ),
    .B(\tcout[2] ),
    .C_N(\tcout[1] ),
    .Y(_098_));
 sky130_fd_sc_hd__nor2_2 _530_ (.A(_336_),
    .B(_382_),
    .Y(_099_));
 sky130_fd_sc_hd__or3_2 _531_ (.A(\tcout[3] ),
    .B(_035_),
    .C(_098_),
    .X(_100_));
 sky130_fd_sc_hd__nand2_2 _532_ (.A(_379_),
    .B(_044_),
    .Y(_101_));
 sky130_fd_sc_hd__a21oi_2 _533_ (.A1(_379_),
    .A2(_044_),
    .B1(_334_),
    .Y(_102_));
 sky130_fd_sc_hd__a221oi_2 _534_ (.A1(_038_),
    .A2(_056_),
    .B1(_100_),
    .B2(_102_),
    .C1(\tcout[5] ),
    .Y(_103_));
 sky130_fd_sc_hd__o211a_2 _535_ (.A1(_018_),
    .A2(_022_),
    .B1(_024_),
    .C1(_376_),
    .X(_104_));
 sky130_fd_sc_hd__or4_2 _536_ (.A(_328_),
    .B(_097_),
    .C(_103_),
    .D(_104_),
    .X(_105_));
 sky130_fd_sc_hd__nor2_2 _537_ (.A(_378_),
    .B(_022_),
    .Y(_106_));
 sky130_fd_sc_hd__a21oi_2 _538_ (.A1(_065_),
    .A2(_089_),
    .B1(_335_),
    .Y(_107_));
 sky130_fd_sc_hd__o21a_2 _539_ (.A1(_106_),
    .A2(_107_),
    .B1(_372_),
    .X(_108_));
 sky130_fd_sc_hd__o211a_2 _540_ (.A1(_335_),
    .A2(_057_),
    .B1(_076_),
    .C1(_362_),
    .X(_109_));
 sky130_fd_sc_hd__o311a_2 _541_ (.A1(_339_),
    .A2(_344_),
    .A3(_382_),
    .B1(_338_),
    .C1(\tcout[4] ),
    .X(_110_));
 sky130_fd_sc_hd__a31o_2 _542_ (.A1(\tcout[3] ),
    .A2(_374_),
    .A3(_381_),
    .B1(_377_),
    .X(_111_));
 sky130_fd_sc_hd__o31ai_2 _543_ (.A1(\tcout[5] ),
    .A2(_109_),
    .A3(_110_),
    .B1(_111_),
    .Y(_112_));
 sky130_fd_sc_hd__o311a_2 _544_ (.A1(\tcout[6] ),
    .A2(_108_),
    .A3(_112_),
    .B1(\tcout[7] ),
    .C1(_105_),
    .X(_113_));
 sky130_fd_sc_hd__a21oi_2 _545_ (.A1(_335_),
    .A2(_019_),
    .B1(_355_),
    .Y(_114_));
 sky130_fd_sc_hd__and3b_2 _546_ (.A_N(\tcout[3] ),
    .B(\tcout[2] ),
    .C(\tcout[1] ),
    .X(_115_));
 sky130_fd_sc_hd__nand3b_2 _547_ (.A_N(\tcout[3] ),
    .B(\tcout[2] ),
    .C(\tcout[1] ),
    .Y(_116_));
 sky130_fd_sc_hd__o311a_2 _548_ (.A1(_366_),
    .A2(_025_),
    .A3(_055_),
    .B1(_116_),
    .C1(\tcout[4] ),
    .X(_117_));
 sky130_fd_sc_hd__o21a_2 _549_ (.A1(_114_),
    .A2(_117_),
    .B1(_333_),
    .X(_118_));
 sky130_fd_sc_hd__o221a_2 _550_ (.A1(\tcout[0] ),
    .A2(_359_),
    .B1(_383_),
    .B2(\tcout[2] ),
    .C1(\tcout[3] ),
    .X(_119_));
 sky130_fd_sc_hd__nor2_2 _551_ (.A(\tcout[3] ),
    .B(_345_),
    .Y(_120_));
 sky130_fd_sc_hd__a21o_2 _552_ (.A1(_374_),
    .A2(_120_),
    .B1(_119_),
    .X(_121_));
 sky130_fd_sc_hd__nand2_2 _553_ (.A(\tcout[2] ),
    .B(_375_),
    .Y(_122_));
 sky130_fd_sc_hd__nand2_2 _554_ (.A(_367_),
    .B(_122_),
    .Y(_123_));
 sky130_fd_sc_hd__a32o_2 _555_ (.A1(_357_),
    .A2(_376_),
    .A3(_123_),
    .B1(_121_),
    .B2(_372_),
    .X(_124_));
 sky130_fd_sc_hd__or3_2 _556_ (.A(_328_),
    .B(_118_),
    .C(_124_),
    .X(_125_));
 sky130_fd_sc_hd__a21o_2 _557_ (.A1(_336_),
    .A2(_375_),
    .B1(_051_),
    .X(_126_));
 sky130_fd_sc_hd__a31o_2 _558_ (.A1(_349_),
    .A2(_381_),
    .A3(_036_),
    .B1(\tcout[3] ),
    .X(_127_));
 sky130_fd_sc_hd__nor2_2 _559_ (.A(_349_),
    .B(_367_),
    .Y(_128_));
 sky130_fd_sc_hd__a21o_2 _560_ (.A1(_126_),
    .A2(_127_),
    .B1(_128_),
    .X(_129_));
 sky130_fd_sc_hd__o221a_2 _561_ (.A1(\tcout[3] ),
    .A2(_019_),
    .B1(_032_),
    .B2(_088_),
    .C1(\tcout[4] ),
    .X(_130_));
 sky130_fd_sc_hd__or3_2 _562_ (.A(\tcout[6] ),
    .B(_333_),
    .C(_130_),
    .X(_131_));
 sky130_fd_sc_hd__o22a_2 _563_ (.A1(_350_),
    .A2(_356_),
    .B1(_375_),
    .B2(_045_),
    .X(_132_));
 sky130_fd_sc_hd__nor2_2 _564_ (.A(\tcout[4] ),
    .B(_132_),
    .Y(_133_));
 sky130_fd_sc_hd__o21ai_2 _565_ (.A1(_366_),
    .A2(_041_),
    .B1(_350_),
    .Y(_134_));
 sky130_fd_sc_hd__a211o_2 _566_ (.A1(_102_),
    .A2(_134_),
    .B1(_133_),
    .C1(_030_),
    .X(_135_));
 sky130_fd_sc_hd__a22o_2 _567_ (.A1(_372_),
    .A2(_129_),
    .B1(_131_),
    .B2(_135_),
    .X(_136_));
 sky130_fd_sc_hd__a31o_2 _568_ (.A1(_337_),
    .A2(_125_),
    .A3(_136_),
    .B1(_113_),
    .X(sine_out[2]));
 sky130_fd_sc_hd__nor3b_2 _569_ (.A(\tcout[0] ),
    .B(\tcout[1] ),
    .C_N(\tcout[2] ),
    .Y(_137_));
 sky130_fd_sc_hd__nor3_2 _570_ (.A(\tcout[3] ),
    .B(_345_),
    .C(_137_),
    .Y(_138_));
 sky130_fd_sc_hd__o21a_2 _571_ (.A1(_119_),
    .A2(_138_),
    .B1(_334_),
    .X(_139_));
 sky130_fd_sc_hd__a21o_2 _572_ (.A1(\tcout[2] ),
    .A2(_001_),
    .B1(\tcout[3] ),
    .X(_140_));
 sky130_fd_sc_hd__or2_2 _573_ (.A(_380_),
    .B(_052_),
    .X(_141_));
 sky130_fd_sc_hd__o211a_2 _574_ (.A1(_035_),
    .A2(_141_),
    .B1(_140_),
    .C1(\tcout[4] ),
    .X(_142_));
 sky130_fd_sc_hd__o21a_2 _575_ (.A1(_139_),
    .A2(_142_),
    .B1(_333_),
    .X(_143_));
 sky130_fd_sc_hd__nand2_2 _576_ (.A(_383_),
    .B(_120_),
    .Y(_144_));
 sky130_fd_sc_hd__a21oi_2 _577_ (.A1(_061_),
    .A2(_144_),
    .B1(_377_),
    .Y(_145_));
 sky130_fd_sc_hd__a211o_2 _578_ (.A1(\tcout[2] ),
    .A2(_001_),
    .B1(_354_),
    .C1(\tcout[3] ),
    .X(_146_));
 sky130_fd_sc_hd__nor2_2 _579_ (.A(_340_),
    .B(_052_),
    .Y(_147_));
 sky130_fd_sc_hd__or3_2 _580_ (.A(_340_),
    .B(_051_),
    .C(_052_),
    .X(_148_));
 sky130_fd_sc_hd__and3_2 _581_ (.A(_372_),
    .B(_146_),
    .C(_148_),
    .X(_149_));
 sky130_fd_sc_hd__or4_2 _582_ (.A(_328_),
    .B(_143_),
    .C(_145_),
    .D(_149_),
    .X(_150_));
 sky130_fd_sc_hd__o21ai_2 _583_ (.A1(_035_),
    .A2(_141_),
    .B1(_362_),
    .Y(_151_));
 sky130_fd_sc_hd__o211a_2 _584_ (.A1(_352_),
    .A2(_032_),
    .B1(_369_),
    .C1(_334_),
    .X(_152_));
 sky130_fd_sc_hd__a211o_2 _585_ (.A1(\tcout[4] ),
    .A2(_151_),
    .B1(_152_),
    .C1(\tcout[5] ),
    .X(_153_));
 sky130_fd_sc_hd__a221o_2 _586_ (.A1(_102_),
    .A2(_134_),
    .B1(_141_),
    .B2(_146_),
    .C1(\tcout[6] ),
    .X(_154_));
 sky130_fd_sc_hd__nand2_2 _587_ (.A(_030_),
    .B(_154_),
    .Y(_155_));
 sky130_fd_sc_hd__a21oi_2 _588_ (.A1(_153_),
    .A2(_155_),
    .B1(\tcout[7] ),
    .Y(_156_));
 sky130_fd_sc_hd__a21oi_2 _589_ (.A1(\tcout[2] ),
    .A2(\tcout[1] ),
    .B1(\tcout[3] ),
    .Y(_157_));
 sky130_fd_sc_hd__nand2_2 _590_ (.A(_089_),
    .B(_157_),
    .Y(_158_));
 sky130_fd_sc_hd__a221o_2 _591_ (.A1(\tcout[4] ),
    .A2(_151_),
    .B1(_158_),
    .B2(_026_),
    .C1(\tcout[5] ),
    .X(_159_));
 sky130_fd_sc_hd__o311a_2 _592_ (.A1(\tcout[4] ),
    .A2(\tcout[1] ),
    .A3(_348_),
    .B1(_045_),
    .C1(\tcout[5] ),
    .X(_160_));
 sky130_fd_sc_hd__nand2_2 _593_ (.A(_134_),
    .B(_160_),
    .Y(_161_));
 sky130_fd_sc_hd__a21o_2 _594_ (.A1(_159_),
    .A2(_161_),
    .B1(\tcout[6] ),
    .X(_162_));
 sky130_fd_sc_hd__o21ai_2 _595_ (.A1(_035_),
    .A2(_052_),
    .B1(_140_),
    .Y(_163_));
 sky130_fd_sc_hd__a21oi_2 _596_ (.A1(_146_),
    .A2(_148_),
    .B1(_373_),
    .Y(_164_));
 sky130_fd_sc_hd__and2_2 _597_ (.A(_339_),
    .B(_353_),
    .X(_165_));
 sky130_fd_sc_hd__nand2_2 _598_ (.A(_339_),
    .B(_001_),
    .Y(_166_));
 sky130_fd_sc_hd__nand2_2 _599_ (.A(_349_),
    .B(_157_),
    .Y(_167_));
 sky130_fd_sc_hd__a31o_2 _600_ (.A1(_046_),
    .A2(_166_),
    .A3(_167_),
    .B1(_377_),
    .X(_168_));
 sky130_fd_sc_hd__or3b_2 _601_ (.A(_328_),
    .B(_164_),
    .C_N(_168_),
    .X(_169_));
 sky130_fd_sc_hd__a31o_2 _602_ (.A1(_333_),
    .A2(_027_),
    .A3(_163_),
    .B1(_169_),
    .X(_170_));
 sky130_fd_sc_hd__a32o_2 _603_ (.A1(\tcout[7] ),
    .A2(_162_),
    .A3(_170_),
    .B1(_150_),
    .B2(_156_),
    .X(sine_out[3]));
 sky130_fd_sc_hd__nor2_2 _604_ (.A(\tcout[4] ),
    .B(_115_),
    .Y(_171_));
 sky130_fd_sc_hd__and3_2 _605_ (.A(_334_),
    .B(_078_),
    .C(_116_),
    .X(_172_));
 sky130_fd_sc_hd__a21o_2 _606_ (.A1(\tcout[2] ),
    .A2(_383_),
    .B1(_368_),
    .X(_173_));
 sky130_fd_sc_hd__a21oi_2 _607_ (.A1(_383_),
    .A2(_044_),
    .B1(_334_),
    .Y(_174_));
 sky130_fd_sc_hd__a22oi_2 _608_ (.A1(_148_),
    .A2(_172_),
    .B1(_173_),
    .B2(_174_),
    .Y(_175_));
 sky130_fd_sc_hd__nor2_2 _609_ (.A(_380_),
    .B(_032_),
    .Y(_176_));
 sky130_fd_sc_hd__o2111a_2 _610_ (.A1(_380_),
    .A2(_032_),
    .B1(\tcout[5] ),
    .C1(_353_),
    .D1(_368_),
    .X(_177_));
 sky130_fd_sc_hd__and3_2 _611_ (.A(\tcout[4] ),
    .B(_353_),
    .C(_361_),
    .X(_178_));
 sky130_fd_sc_hd__o31ai_2 _612_ (.A1(\tcout[0] ),
    .A2(\tcout[2] ),
    .A3(\tcout[1] ),
    .B1(\tcout[3] ),
    .Y(_179_));
 sky130_fd_sc_hd__a2bb2o_2 _613_ (.A1_N(_376_),
    .A2_N(_177_),
    .B1(_178_),
    .B2(_179_),
    .X(_180_));
 sky130_fd_sc_hd__o211a_2 _614_ (.A1(\tcout[5] ),
    .A2(_175_),
    .B1(_180_),
    .C1(\tcout[6] ),
    .X(_181_));
 sky130_fd_sc_hd__o211a_2 _615_ (.A1(\tcout[2] ),
    .A2(_001_),
    .B1(_050_),
    .C1(_335_),
    .X(_182_));
 sky130_fd_sc_hd__a211o_2 _616_ (.A1(_122_),
    .A2(_147_),
    .B1(_182_),
    .C1(_373_),
    .X(_183_));
 sky130_fd_sc_hd__o211ai_2 _617_ (.A1(\tcout[2] ),
    .A2(_375_),
    .B1(_359_),
    .C1(\tcout[3] ),
    .Y(_184_));
 sky130_fd_sc_hd__a31o_2 _618_ (.A1(_367_),
    .A2(_042_),
    .A3(_184_),
    .B1(_377_),
    .X(_185_));
 sky130_fd_sc_hd__and3_2 _619_ (.A(_328_),
    .B(_183_),
    .C(_185_),
    .X(_186_));
 sky130_fd_sc_hd__nand4_2 _620_ (.A(_338_),
    .B(_032_),
    .C(_066_),
    .D(_078_),
    .Y(_187_));
 sky130_fd_sc_hd__a31o_2 _621_ (.A1(\tcout[3] ),
    .A2(_346_),
    .A3(_361_),
    .B1(\tcout[4] ),
    .X(_188_));
 sky130_fd_sc_hd__a21o_2 _622_ (.A1(_187_),
    .A2(_188_),
    .B1(\tcout[5] ),
    .X(_189_));
 sky130_fd_sc_hd__a21oi_2 _623_ (.A1(_186_),
    .A2(_189_),
    .B1(_181_),
    .Y(_190_));
 sky130_fd_sc_hd__a31o_2 _624_ (.A1(_346_),
    .A2(_361_),
    .A3(_367_),
    .B1(\tcout[4] ),
    .X(_191_));
 sky130_fd_sc_hd__a21o_2 _625_ (.A1(_187_),
    .A2(_191_),
    .B1(_030_),
    .X(_192_));
 sky130_fd_sc_hd__o211a_2 _626_ (.A1(_181_),
    .A2(_186_),
    .B1(_192_),
    .C1(\tcout[7] ),
    .X(_193_));
 sky130_fd_sc_hd__a21oi_2 _627_ (.A1(_337_),
    .A2(_190_),
    .B1(_193_),
    .Y(sine_out[4]));
 sky130_fd_sc_hd__o211ai_2 _628_ (.A1(_021_),
    .A2(_032_),
    .B1(_134_),
    .C1(\tcout[4] ),
    .Y(_194_));
 sky130_fd_sc_hd__nand2_2 _629_ (.A(_076_),
    .B(_184_),
    .Y(_195_));
 sky130_fd_sc_hd__a21oi_2 _630_ (.A1(_194_),
    .A2(_195_),
    .B1(_030_),
    .Y(_196_));
 sky130_fd_sc_hd__and4_2 _631_ (.A(_335_),
    .B(_349_),
    .C(_381_),
    .D(_036_),
    .X(_197_));
 sky130_fd_sc_hd__nand2_2 _632_ (.A(_028_),
    .B(_102_),
    .Y(_198_));
 sky130_fd_sc_hd__nor2_2 _633_ (.A(\tcout[6] ),
    .B(_373_),
    .Y(_199_));
 sky130_fd_sc_hd__or4b_2 _634_ (.A(_055_),
    .B(_137_),
    .C(_176_),
    .D_N(_199_),
    .X(_200_));
 sky130_fd_sc_hd__o21ai_2 _635_ (.A1(_197_),
    .A2(_198_),
    .B1(_200_),
    .Y(_201_));
 sky130_fd_sc_hd__a32o_2 _636_ (.A1(\tcout[3] ),
    .A2(_089_),
    .A3(_122_),
    .B1(_120_),
    .B2(_374_),
    .X(_202_));
 sky130_fd_sc_hd__o211a_2 _637_ (.A1(_349_),
    .A2(_367_),
    .B1(\tcout[4] ),
    .C1(_338_),
    .X(_203_));
 sky130_fd_sc_hd__a31o_2 _638_ (.A1(_370_),
    .A2(_122_),
    .A3(_203_),
    .B1(\tcout[5] ),
    .X(_204_));
 sky130_fd_sc_hd__a21o_2 _639_ (.A1(_334_),
    .A2(_202_),
    .B1(_204_),
    .X(_205_));
 sky130_fd_sc_hd__and2_2 _640_ (.A(_343_),
    .B(_370_),
    .X(_206_));
 sky130_fd_sc_hd__nand2_2 _641_ (.A(\tcout[0] ),
    .B(_342_),
    .Y(_207_));
 sky130_fd_sc_hd__o2111a_2 _642_ (.A1(_339_),
    .A2(_379_),
    .B1(_207_),
    .C1(_357_),
    .D1(_334_),
    .X(_208_));
 sky130_fd_sc_hd__a311o_2 _643_ (.A1(\tcout[4] ),
    .A2(_158_),
    .A3(_206_),
    .B1(_208_),
    .C1(_333_),
    .X(_209_));
 sky130_fd_sc_hd__a31o_2 _644_ (.A1(\tcout[6] ),
    .A2(_205_),
    .A3(_209_),
    .B1(_201_),
    .X(_210_));
 sky130_fd_sc_hd__a311o_2 _645_ (.A1(\tcout[6] ),
    .A2(_205_),
    .A3(_209_),
    .B1(_196_),
    .C1(_201_),
    .X(_211_));
 sky130_fd_sc_hd__a31o_2 _646_ (.A1(_046_),
    .A2(_086_),
    .A3(_166_),
    .B1(\tcout[4] ),
    .X(_212_));
 sky130_fd_sc_hd__a21o_2 _647_ (.A1(_194_),
    .A2(_212_),
    .B1(_030_),
    .X(_213_));
 sky130_fd_sc_hd__nand2_2 _648_ (.A(\tcout[7] ),
    .B(_213_),
    .Y(_214_));
 sky130_fd_sc_hd__o2bb2a_2 _649_ (.A1_N(_337_),
    .A2_N(_211_),
    .B1(_214_),
    .B2(_210_),
    .X(sine_out[5]));
 sky130_fd_sc_hd__a221o_2 _650_ (.A1(_352_),
    .A2(_041_),
    .B1(_051_),
    .B2(_335_),
    .C1(\tcout[4] ),
    .X(_215_));
 sky130_fd_sc_hd__a31oi_2 _651_ (.A1(\tcout[3] ),
    .A2(_346_),
    .A3(_122_),
    .B1(_215_),
    .Y(_216_));
 sky130_fd_sc_hd__nand2_2 _652_ (.A(_001_),
    .B(_041_),
    .Y(_217_));
 sky130_fd_sc_hd__a41o_2 _653_ (.A1(\tcout[4] ),
    .A2(_365_),
    .A3(_207_),
    .A4(_217_),
    .B1(\tcout[5] ),
    .X(_218_));
 sky130_fd_sc_hd__nor2_2 _654_ (.A(_340_),
    .B(_001_),
    .Y(_219_));
 sky130_fd_sc_hd__nor2_2 _655_ (.A(\tcout[3] ),
    .B(_021_),
    .Y(_220_));
 sky130_fd_sc_hd__o21ai_2 _656_ (.A1(_219_),
    .A2(_220_),
    .B1(_376_),
    .Y(_221_));
 sky130_fd_sc_hd__a21oi_2 _657_ (.A1(_089_),
    .A2(_122_),
    .B1(_335_),
    .Y(_222_));
 sky130_fd_sc_hd__o211ai_2 _658_ (.A1(_335_),
    .A2(_122_),
    .B1(_089_),
    .C1(_372_),
    .Y(_223_));
 sky130_fd_sc_hd__o211ai_2 _659_ (.A1(_216_),
    .A2(_218_),
    .B1(_221_),
    .C1(_223_),
    .Y(_224_));
 sky130_fd_sc_hd__o211a_2 _660_ (.A1(\tcout[2] ),
    .A2(_383_),
    .B1(_359_),
    .C1(\tcout[3] ),
    .X(_225_));
 sky130_fd_sc_hd__or3b_2 _661_ (.A(_373_),
    .B(_225_),
    .C_N(_369_),
    .X(_226_));
 sky130_fd_sc_hd__a211o_2 _662_ (.A1(_383_),
    .A2(_044_),
    .B1(_358_),
    .C1(_377_),
    .X(_227_));
 sky130_fd_sc_hd__a21oi_2 _663_ (.A1(_226_),
    .A2(_227_),
    .B1(\tcout[6] ),
    .Y(_228_));
 sky130_fd_sc_hd__a21o_2 _664_ (.A1(_049_),
    .A2(_173_),
    .B1(_334_),
    .X(_229_));
 sky130_fd_sc_hd__a21o_2 _665_ (.A1(_356_),
    .A2(_179_),
    .B1(\tcout[4] ),
    .X(_230_));
 sky130_fd_sc_hd__a21oi_2 _666_ (.A1(_229_),
    .A2(_230_),
    .B1(_030_),
    .Y(_231_));
 sky130_fd_sc_hd__a211oi_2 _667_ (.A1(\tcout[6] ),
    .A2(_224_),
    .B1(_228_),
    .C1(_231_),
    .Y(_232_));
 sky130_fd_sc_hd__o31ai_2 _668_ (.A1(\tcout[4] ),
    .A2(_366_),
    .A3(_021_),
    .B1(_229_),
    .Y(_233_));
 sky130_fd_sc_hd__a221o_2 _669_ (.A1(\tcout[6] ),
    .A2(_224_),
    .B1(_233_),
    .B2(_029_),
    .C1(_228_),
    .X(_234_));
 sky130_fd_sc_hd__mux2_1 _670_ (.A0(_232_),
    .A1(_234_),
    .S(\tcout[7] ),
    .X(sine_out[6]));
 sky130_fd_sc_hd__a31o_2 _671_ (.A1(_335_),
    .A2(\tcout[2] ),
    .A3(_379_),
    .B1(\tcout[4] ),
    .X(_235_));
 sky130_fd_sc_hd__o32a_2 _672_ (.A1(_334_),
    .A2(_021_),
    .A3(_055_),
    .B1(_096_),
    .B2(_235_),
    .X(_236_));
 sky130_fd_sc_hd__o31ai_2 _673_ (.A1(_377_),
    .A2(_051_),
    .A3(_220_),
    .B1(\tcout[6] ),
    .Y(_237_));
 sky130_fd_sc_hd__a21oi_2 _674_ (.A1(_336_),
    .A2(_383_),
    .B1(_022_),
    .Y(_238_));
 sky130_fd_sc_hd__a21o_2 _675_ (.A1(_379_),
    .A2(_031_),
    .B1(_373_),
    .X(_239_));
 sky130_fd_sc_hd__o22ai_2 _676_ (.A1(\tcout[5] ),
    .A2(_236_),
    .B1(_238_),
    .B2(_239_),
    .Y(_240_));
 sky130_fd_sc_hd__a2111o_2 _677_ (.A1(\tcout[1] ),
    .A2(_344_),
    .B1(_345_),
    .C1(_382_),
    .D1(_335_),
    .X(_241_));
 sky130_fd_sc_hd__a32o_2 _678_ (.A1(_334_),
    .A2(_042_),
    .A3(_179_),
    .B1(_241_),
    .B2(_066_),
    .X(_242_));
 sky130_fd_sc_hd__and2_2 _679_ (.A(_333_),
    .B(_242_),
    .X(_243_));
 sky130_fd_sc_hd__or3_2 _680_ (.A(\tcout[3] ),
    .B(_352_),
    .C(_380_),
    .X(_244_));
 sky130_fd_sc_hd__o21a_2 _681_ (.A1(_051_),
    .A2(_052_),
    .B1(_376_),
    .X(_245_));
 sky130_fd_sc_hd__a221o_2 _682_ (.A1(_372_),
    .A2(_206_),
    .B1(_244_),
    .B2(_245_),
    .C1(\tcout[6] ),
    .X(_246_));
 sky130_fd_sc_hd__o22a_2 _683_ (.A1(_237_),
    .A2(_240_),
    .B1(_243_),
    .B2(_246_),
    .X(_247_));
 sky130_fd_sc_hd__nand2_2 _684_ (.A(_021_),
    .B(_038_),
    .Y(_248_));
 sky130_fd_sc_hd__and2_2 _685_ (.A(\tcout[7] ),
    .B(_248_),
    .X(_249_));
 sky130_fd_sc_hd__mux2_1 _686_ (.A0(_249_),
    .A1(_337_),
    .S(_247_),
    .X(sine_out[7]));
 sky130_fd_sc_hd__o21ai_2 _687_ (.A1(\tcout[4] ),
    .A2(_023_),
    .B1(_028_),
    .Y(_250_));
 sky130_fd_sc_hd__a31o_2 _688_ (.A1(\tcout[4] ),
    .A2(_144_),
    .A3(_166_),
    .B1(_250_),
    .X(_251_));
 sky130_fd_sc_hd__a22o_2 _689_ (.A1(\tcout[4] ),
    .A2(_062_),
    .B1(_079_),
    .B2(_171_),
    .X(_252_));
 sky130_fd_sc_hd__o21a_2 _690_ (.A1(\tcout[0] ),
    .A2(_368_),
    .B1(_370_),
    .X(_253_));
 sky130_fd_sc_hd__o21ai_2 _691_ (.A1(_377_),
    .A2(_253_),
    .B1(\tcout[6] ),
    .Y(_254_));
 sky130_fd_sc_hd__or3_2 _692_ (.A(_335_),
    .B(_350_),
    .C(_352_),
    .X(_255_));
 sky130_fd_sc_hd__o211a_2 _693_ (.A1(_137_),
    .A2(_244_),
    .B1(_255_),
    .C1(_372_),
    .X(_256_));
 sky130_fd_sc_hd__a211o_2 _694_ (.A1(_333_),
    .A2(_252_),
    .B1(_254_),
    .C1(_256_),
    .X(_257_));
 sky130_fd_sc_hd__nand2_2 _695_ (.A(_251_),
    .B(_257_),
    .Y(_258_));
 sky130_fd_sc_hd__o21ai_2 _696_ (.A1(\tcout[3] ),
    .A2(_374_),
    .B1(_381_),
    .Y(_259_));
 sky130_fd_sc_hd__o221a_2 _697_ (.A1(_346_),
    .A2(_367_),
    .B1(_259_),
    .B2(_352_),
    .C1(\tcout[4] ),
    .X(_260_));
 sky130_fd_sc_hd__a21oi_2 _698_ (.A1(_086_),
    .A2(_206_),
    .B1(\tcout[4] ),
    .Y(_261_));
 sky130_fd_sc_hd__o21a_2 _699_ (.A1(_260_),
    .A2(_261_),
    .B1(_029_),
    .X(_262_));
 sky130_fd_sc_hd__o21a_2 _700_ (.A1(\tcout[0] ),
    .A2(_095_),
    .B1(_076_),
    .X(_263_));
 sky130_fd_sc_hd__o21ai_2 _701_ (.A1(_260_),
    .A2(_263_),
    .B1(_029_),
    .Y(_264_));
 sky130_fd_sc_hd__a31o_2 _702_ (.A1(_251_),
    .A2(_257_),
    .A3(_264_),
    .B1(\tcout[7] ),
    .X(_265_));
 sky130_fd_sc_hd__o31a_2 _703_ (.A1(_337_),
    .A2(_258_),
    .A3(_262_),
    .B1(_265_),
    .X(sine_out[8]));
 sky130_fd_sc_hd__a21o_2 _704_ (.A1(\tcout[0] ),
    .A2(\tcout[3] ),
    .B1(_197_),
    .X(_266_));
 sky130_fd_sc_hd__o211a_2 _705_ (.A1(_340_),
    .A2(_001_),
    .B1(_334_),
    .C1(\tcout[3] ),
    .X(_267_));
 sky130_fd_sc_hd__a211o_2 _706_ (.A1(\tcout[4] ),
    .A2(_266_),
    .B1(_267_),
    .C1(\tcout[5] ),
    .X(_268_));
 sky130_fd_sc_hd__a21o_2 _707_ (.A1(_023_),
    .A2(_063_),
    .B1(_377_),
    .X(_269_));
 sky130_fd_sc_hd__o22a_2 _708_ (.A1(_335_),
    .A2(_050_),
    .B1(_088_),
    .B2(_099_),
    .X(_270_));
 sky130_fd_sc_hd__o311a_2 _709_ (.A1(_373_),
    .A2(_054_),
    .A3(_270_),
    .B1(_269_),
    .C1(\tcout[6] ),
    .X(_271_));
 sky130_fd_sc_hd__a21oi_2 _710_ (.A1(_356_),
    .A2(_179_),
    .B1(_377_),
    .Y(_272_));
 sky130_fd_sc_hd__nor2_2 _711_ (.A(\tcout[6] ),
    .B(_272_),
    .Y(_273_));
 sky130_fd_sc_hd__o311a_2 _712_ (.A1(_041_),
    .A2(_088_),
    .A3(_099_),
    .B1(_217_),
    .C1(\tcout[4] ),
    .X(_274_));
 sky130_fd_sc_hd__a31o_2 _713_ (.A1(_334_),
    .A2(_023_),
    .A3(_063_),
    .B1(\tcout[5] ),
    .X(_275_));
 sky130_fd_sc_hd__o32a_2 _714_ (.A1(_373_),
    .A2(_055_),
    .A3(_222_),
    .B1(_274_),
    .B2(_275_),
    .X(_276_));
 sky130_fd_sc_hd__a22o_2 _715_ (.A1(_268_),
    .A2(_271_),
    .B1(_273_),
    .B2(_276_),
    .X(_277_));
 sky130_fd_sc_hd__mux2_1 _716_ (.A0(_337_),
    .A1(_249_),
    .S(_277_),
    .X(sine_out[9]));
 sky130_fd_sc_hd__or2_2 _717_ (.A(_354_),
    .B(_057_),
    .X(_002_));
 sky130_fd_sc_hd__o211a_2 _718_ (.A1(_018_),
    .A2(_022_),
    .B1(\tcout[4] ),
    .C1(_338_),
    .X(_278_));
 sky130_fd_sc_hd__o31ai_2 _719_ (.A1(\tcout[4] ),
    .A2(_354_),
    .A3(_057_),
    .B1(_333_),
    .Y(_279_));
 sky130_fd_sc_hd__a21o_2 _720_ (.A1(_351_),
    .A2(_127_),
    .B1(_377_),
    .X(_280_));
 sky130_fd_sc_hd__a31o_2 _721_ (.A1(_341_),
    .A2(_001_),
    .A3(_049_),
    .B1(_239_),
    .X(_281_));
 sky130_fd_sc_hd__o31a_2 _722_ (.A1(_038_),
    .A2(_278_),
    .A3(_279_),
    .B1(\tcout[6] ),
    .X(_282_));
 sky130_fd_sc_hd__nor2_2 _723_ (.A(_057_),
    .B(_179_),
    .Y(_283_));
 sky130_fd_sc_hd__or3_2 _724_ (.A(\tcout[3] ),
    .B(_377_),
    .C(_018_),
    .X(_284_));
 sky130_fd_sc_hd__o311a_2 _725_ (.A1(_373_),
    .A2(_062_),
    .A3(_283_),
    .B1(_284_),
    .C1(_328_),
    .X(_285_));
 sky130_fd_sc_hd__a31o_2 _726_ (.A1(_280_),
    .A2(_281_),
    .A3(_282_),
    .B1(_285_),
    .X(_286_));
 sky130_fd_sc_hd__a22o_2 _727_ (.A1(\tcout[2] ),
    .A2(_379_),
    .B1(_383_),
    .B2(\tcout[3] ),
    .X(_287_));
 sky130_fd_sc_hd__a211o_2 _728_ (.A1(_101_),
    .A2(_287_),
    .B1(_334_),
    .C1(_098_),
    .X(_288_));
 sky130_fd_sc_hd__a31o_2 _729_ (.A1(\tcout[3] ),
    .A2(_089_),
    .A3(_122_),
    .B1(_081_),
    .X(_289_));
 sky130_fd_sc_hd__nand2_2 _730_ (.A(_334_),
    .B(_289_),
    .Y(_290_));
 sky130_fd_sc_hd__a21oi_2 _731_ (.A1(_288_),
    .A2(_290_),
    .B1(_030_),
    .Y(_291_));
 sky130_fd_sc_hd__nand2_2 _732_ (.A(\tcout[7] ),
    .B(_286_),
    .Y(_292_));
 sky130_fd_sc_hd__o31a_2 _733_ (.A1(_128_),
    .A2(_222_),
    .A3(_235_),
    .B1(_288_),
    .X(_293_));
 sky130_fd_sc_hd__o21a_2 _734_ (.A1(_030_),
    .A2(_293_),
    .B1(_286_),
    .X(_294_));
 sky130_fd_sc_hd__o22a_2 _735_ (.A1(_291_),
    .A2(_292_),
    .B1(_294_),
    .B2(\tcout[7] ),
    .X(sine_out[10]));
 sky130_fd_sc_hd__or3_2 _736_ (.A(\tcout[3] ),
    .B(_360_),
    .C(_021_),
    .X(_295_));
 sky130_fd_sc_hd__a21o_2 _737_ (.A1(_184_),
    .A2(_295_),
    .B1(_377_),
    .X(_296_));
 sky130_fd_sc_hd__o32a_2 _738_ (.A1(_335_),
    .A2(_345_),
    .A3(_360_),
    .B1(_018_),
    .B2(_022_),
    .X(_297_));
 sky130_fd_sc_hd__or3b_2 _739_ (.A(_342_),
    .B(_373_),
    .C_N(_297_),
    .X(_298_));
 sky130_fd_sc_hd__o21a_2 _740_ (.A1(_018_),
    .A2(_055_),
    .B1(_042_),
    .X(_299_));
 sky130_fd_sc_hd__o31a_2 _741_ (.A1(\tcout[4] ),
    .A2(_347_),
    .A3(_023_),
    .B1(_333_),
    .X(_300_));
 sky130_fd_sc_hd__o21ai_2 _742_ (.A1(_334_),
    .A2(_299_),
    .B1(_300_),
    .Y(_301_));
 sky130_fd_sc_hd__a31oi_2 _743_ (.A1(_296_),
    .A2(_298_),
    .A3(_301_),
    .B1(_328_),
    .Y(_302_));
 sky130_fd_sc_hd__a21oi_2 _744_ (.A1(_335_),
    .A2(_002_),
    .B1(_044_),
    .Y(_303_));
 sky130_fd_sc_hd__or4_2 _745_ (.A(_334_),
    .B(\tcout[3] ),
    .C(\tcout[2] ),
    .D(\tcout[1] ),
    .X(_304_));
 sky130_fd_sc_hd__o211a_2 _746_ (.A1(\tcout[4] ),
    .A2(_303_),
    .B1(_304_),
    .C1(_028_),
    .X(_305_));
 sky130_fd_sc_hd__a31o_2 _747_ (.A1(_341_),
    .A2(_349_),
    .A3(_157_),
    .B1(_283_),
    .X(_306_));
 sky130_fd_sc_hd__a22o_2 _748_ (.A1(_148_),
    .A2(_172_),
    .B1(_306_),
    .B2(\tcout[4] ),
    .X(_307_));
 sky130_fd_sc_hd__a211o_2 _749_ (.A1(_029_),
    .A2(_307_),
    .B1(_305_),
    .C1(_302_),
    .X(_308_));
 sky130_fd_sc_hd__mux2_1 _750_ (.A0(_249_),
    .A1(_337_),
    .S(_308_),
    .X(sine_out[11]));
 sky130_fd_sc_hd__mux2_1 _751_ (.A0(_359_),
    .A1(_051_),
    .S(_335_),
    .X(_309_));
 sky130_fd_sc_hd__a21o_2 _752_ (.A1(\tcout[4] ),
    .A2(_309_),
    .B1(\tcout[5] ),
    .X(_310_));
 sky130_fd_sc_hd__a211o_2 _753_ (.A1(_335_),
    .A2(_051_),
    .B1(_165_),
    .C1(\tcout[4] ),
    .X(_311_));
 sky130_fd_sc_hd__a32o_2 _754_ (.A1(_335_),
    .A2(_346_),
    .A3(_018_),
    .B1(_353_),
    .B2(_339_),
    .X(_312_));
 sky130_fd_sc_hd__a21oi_2 _755_ (.A1(_376_),
    .A2(_312_),
    .B1(_328_),
    .Y(_313_));
 sky130_fd_sc_hd__and3_2 _756_ (.A(_310_),
    .B(_311_),
    .C(_313_),
    .X(_314_));
 sky130_fd_sc_hd__o21ai_2 _757_ (.A1(_115_),
    .A2(_165_),
    .B1(_334_),
    .Y(_315_));
 sky130_fd_sc_hd__o311a_2 _758_ (.A1(_334_),
    .A2(_339_),
    .A3(_115_),
    .B1(_315_),
    .C1(_029_),
    .X(_316_));
 sky130_fd_sc_hd__a311o_2 _759_ (.A1(_045_),
    .A2(_078_),
    .A3(_199_),
    .B1(_314_),
    .C1(_316_),
    .X(_317_));
 sky130_fd_sc_hd__a21oi_2 _760_ (.A1(_335_),
    .A2(_021_),
    .B1(_337_),
    .Y(_318_));
 sky130_fd_sc_hd__mux2_1 _761_ (.A0(_337_),
    .A1(_318_),
    .S(_317_),
    .X(sine_out[12]));
 sky130_fd_sc_hd__or2_2 _762_ (.A(_334_),
    .B(_157_),
    .X(_319_));
 sky130_fd_sc_hd__or2_2 _763_ (.A(\tcout[4] ),
    .B(_147_),
    .X(_320_));
 sky130_fd_sc_hd__a221o_2 _764_ (.A1(_333_),
    .A2(_046_),
    .B1(_319_),
    .B2(_320_),
    .C1(_328_),
    .X(_321_));
 sky130_fd_sc_hd__o21ai_2 _765_ (.A1(_165_),
    .A2(_220_),
    .B1(_334_),
    .Y(_322_));
 sky130_fd_sc_hd__a21o_2 _766_ (.A1(_319_),
    .A2(_322_),
    .B1(_030_),
    .X(_323_));
 sky130_fd_sc_hd__o311a_2 _767_ (.A1(\tcout[6] ),
    .A2(_373_),
    .A3(_078_),
    .B1(_321_),
    .C1(_323_),
    .X(_324_));
 sky130_fd_sc_hd__o21a_2 _768_ (.A1(_030_),
    .A2(_248_),
    .B1(_337_),
    .X(_325_));
 sky130_fd_sc_hd__mux2_1 _769_ (.A0(\tcout[7] ),
    .A1(_325_),
    .S(_324_),
    .X(sine_out[13]));
 sky130_fd_sc_hd__o211a_2 _770_ (.A1(\tcout[4] ),
    .A2(_147_),
    .B1(\tcout[6] ),
    .C1(\tcout[5] ),
    .X(_326_));
 sky130_fd_sc_hd__a31o_2 _771_ (.A1(_029_),
    .A2(_248_),
    .A3(_319_),
    .B1(_326_),
    .X(_327_));
 sky130_fd_sc_hd__mux2_1 _772_ (.A0(_325_),
    .A1(\tcout[7] ),
    .S(_327_),
    .X(sine_out[14]));
 sky130_fd_sc_hd__o21a_2 _773_ (.A1(_030_),
    .A2(_248_),
    .B1(\tcout[7] ),
    .X(sine_out[15]));
 sky130_fd_sc_hd__o211ai_2 _774_ (.A1(_347_),
    .A2(_367_),
    .B1(_032_),
    .C1(_338_),
    .Y(_003_));
 sky130_fd_sc_hd__and3_2 _775_ (.A(\tcout[4] ),
    .B(_352_),
    .C(_044_),
    .X(_329_));
 sky130_fd_sc_hd__a21o_2 _776_ (.A1(_352_),
    .A2(_044_),
    .B1(\tcout[4] ),
    .X(_330_));
 sky130_fd_sc_hd__and2b_2 _777_ (.A_N(_329_),
    .B(_330_),
    .X(_004_));
 sky130_fd_sc_hd__xnor2_2 _778_ (.A(_333_),
    .B(_329_),
    .Y(_005_));
 sky130_fd_sc_hd__and3_2 _779_ (.A(\tcout[6] ),
    .B(\tcout[5] ),
    .C(_329_),
    .X(_331_));
 sky130_fd_sc_hd__a21oi_2 _780_ (.A1(\tcout[5] ),
    .A2(_329_),
    .B1(\tcout[6] ),
    .Y(_332_));
 sky130_fd_sc_hd__nor2_2 _781_ (.A(_331_),
    .B(_332_),
    .Y(_006_));
 sky130_fd_sc_hd__xnor2_2 _782_ (.A(_337_),
    .B(_331_),
    .Y(_007_));
 sky130_fd_sc_hd__inv_2 _783_ (.A(rst),
    .Y(_009_));
 sky130_fd_sc_hd__inv_2 _784_ (.A(rst),
    .Y(_010_));
 sky130_fd_sc_hd__inv_2 _785_ (.A(rst),
    .Y(_011_));
 sky130_fd_sc_hd__inv_2 _786_ (.A(rst),
    .Y(_012_));
 sky130_fd_sc_hd__inv_2 _787_ (.A(rst),
    .Y(_013_));
 sky130_fd_sc_hd__inv_2 _788_ (.A(rst),
    .Y(_014_));
 sky130_fd_sc_hd__inv_2 _789_ (.A(rst),
    .Y(_015_));
 sky130_fd_sc_hd__dfrtp_2 _790_ (.CLK(clk),
    .D(_000_),
    .RESET_B(_008_),
    .Q(\tcout[0] ));
 sky130_fd_sc_hd__dfrtp_2 _791_ (.CLK(clk),
    .D(_001_),
    .RESET_B(_009_),
    .Q(\tcout[1] ));
 sky130_fd_sc_hd__dfrtp_2 _792_ (.CLK(clk),
    .D(_002_),
    .RESET_B(_010_),
    .Q(\tcout[2] ));
 sky130_fd_sc_hd__dfrtp_2 _793_ (.CLK(clk),
    .D(_003_),
    .RESET_B(_011_),
    .Q(\tcout[3] ));
 sky130_fd_sc_hd__dfrtp_2 _794_ (.CLK(clk),
    .D(_004_),
    .RESET_B(_012_),
    .Q(\tcout[4] ));
 sky130_fd_sc_hd__dfrtp_2 _795_ (.CLK(clk),
    .D(_005_),
    .RESET_B(_013_),
    .Q(\tcout[5] ));
 sky130_fd_sc_hd__dfrtp_2 _796_ (.CLK(clk),
    .D(_006_),
    .RESET_B(_014_),
    .Q(\tcout[6] ));
 sky130_fd_sc_hd__dfrtp_2 _797_ (.CLK(clk),
    .D(_007_),
    .RESET_B(_015_),
    .Q(\tcout[7] ));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_160 ();
endmodule
